* NGSPICE file created from life_cell.ext - technology: sky130A

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.312 ps=1.62 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203 ps=1.27 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt life_cell VGND VPWR clk d dl dr in_data l load_in load_out out_data prev_out_data
+ r reset run shift state u ul ur vccd1 vssd1
XFILLER_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_49_ net17 net5 VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__nor2_1
XFILLER_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_65_ clknet_1_0__leaf_clk _01_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_48_ _12_ _17_ VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__nand2_1
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_64_ clknet_1_1__leaf_clk _00_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_47_ _14_ _16_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_63_ net7 _30_ _31_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__o21a_1
XFILLER_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_46_ _04_ _08_ _15_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__o21a_1
XFILLER_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_62_ _24_ net7 net10 VGND VGND VPWR VPWR _31_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_45_ _05_ _07_ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__or2_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_61_ net16 net8 net12 VGND VGND VPWR VPWR _30_ sky130_fd_sc_hd__mux2_1
XFILLER_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_44_ net9 _06_ _13_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_60_ _27_ _29_ net10 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_43_ net1 net13 VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__and2_1
XFILLER_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_42_ _02_ _10_ _11_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__o21a_1
XFILLER_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR out_data sky130_fd_sc_hd__buf_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_41_ _03_ _09_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__or2_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput17 net17 VGND VGND VPWR VPWR state sky130_fd_sc_hd__buf_2
XFILLER_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_40_ _03_ _09_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 d VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 dl VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 dr VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 in_data VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 l VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_59_ net11 _28_ VGND VGND VPWR VPWR _29_ sky130_fd_sc_hd__or2b_1
XFILLER_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 load_in VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_58_ net17 net4 net6 VGND VGND VPWR VPWR _28_ sky130_fd_sc_hd__mux2_1
XFILLER_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 load_out VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_57_ _18_ _21_ _23_ _26_ VGND VGND VPWR VPWR _27_ sky130_fd_sc_hd__a211o_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 reset VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 prev_out_data VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_56_ _24_ _25_ _20_ _17_ _12_ VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__o311a_1
XFILLER_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_39_ _04_ _08_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__xnor2_1
Xinput11 run VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 r VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_55_ net5 VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__inv_2
XFILLER_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 shift VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
XFILLER_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_38_ _05_ _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_54_ net17 VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__inv_2
XFILLER_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 u VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_37_ net9 _06_ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_53_ _12_ _17_ _22_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 ul VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_36_ net1 net13 VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__xor2_1
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ _14_ _16_ net11 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__o21a_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput15 ur VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_35_ net2 VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__inv_2
XFILLER_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_51_ net5 _19_ _20_ VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__mux2_1
XFILLER_23_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34_ net15 VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__inv_2
XFILLER_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_50_ _02_ _10_ VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_33_ net14 VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__inv_2
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_32_ net3 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__inv_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
.ends

