module game_of_life (clk,
    inp_load,
    out_load,
    out_shift,
    reset,
    run,
    inp_data,
    inp_y_addr,
    out_data);
 input clk;
 input inp_load;
 input out_load;
 input out_shift;
 input reset;
 input run;
 input [15:0] inp_data;
 input [3:0] inp_y_addr;
 output [15:0] out_data;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire \cell_outs[0] ;
 wire \cell_outs[100] ;
 wire \cell_outs[101] ;
 wire \cell_outs[102] ;
 wire \cell_outs[103] ;
 wire \cell_outs[104] ;
 wire \cell_outs[105] ;
 wire \cell_outs[106] ;
 wire \cell_outs[107] ;
 wire \cell_outs[108] ;
 wire \cell_outs[109] ;
 wire \cell_outs[10] ;
 wire \cell_outs[110] ;
 wire \cell_outs[111] ;
 wire \cell_outs[112] ;
 wire \cell_outs[113] ;
 wire \cell_outs[114] ;
 wire \cell_outs[115] ;
 wire \cell_outs[116] ;
 wire \cell_outs[117] ;
 wire \cell_outs[118] ;
 wire \cell_outs[119] ;
 wire \cell_outs[11] ;
 wire \cell_outs[120] ;
 wire \cell_outs[121] ;
 wire \cell_outs[122] ;
 wire \cell_outs[123] ;
 wire \cell_outs[124] ;
 wire \cell_outs[125] ;
 wire \cell_outs[126] ;
 wire \cell_outs[127] ;
 wire \cell_outs[128] ;
 wire \cell_outs[129] ;
 wire \cell_outs[12] ;
 wire \cell_outs[130] ;
 wire \cell_outs[131] ;
 wire \cell_outs[132] ;
 wire \cell_outs[133] ;
 wire \cell_outs[134] ;
 wire \cell_outs[135] ;
 wire \cell_outs[136] ;
 wire \cell_outs[137] ;
 wire \cell_outs[138] ;
 wire \cell_outs[139] ;
 wire \cell_outs[13] ;
 wire \cell_outs[140] ;
 wire \cell_outs[141] ;
 wire \cell_outs[142] ;
 wire \cell_outs[143] ;
 wire \cell_outs[144] ;
 wire \cell_outs[145] ;
 wire \cell_outs[146] ;
 wire \cell_outs[147] ;
 wire \cell_outs[148] ;
 wire \cell_outs[149] ;
 wire \cell_outs[14] ;
 wire \cell_outs[150] ;
 wire \cell_outs[151] ;
 wire \cell_outs[152] ;
 wire \cell_outs[153] ;
 wire \cell_outs[154] ;
 wire \cell_outs[155] ;
 wire \cell_outs[156] ;
 wire \cell_outs[157] ;
 wire \cell_outs[158] ;
 wire \cell_outs[159] ;
 wire \cell_outs[15] ;
 wire \cell_outs[160] ;
 wire \cell_outs[161] ;
 wire \cell_outs[162] ;
 wire \cell_outs[163] ;
 wire \cell_outs[164] ;
 wire \cell_outs[165] ;
 wire \cell_outs[166] ;
 wire \cell_outs[167] ;
 wire \cell_outs[168] ;
 wire \cell_outs[169] ;
 wire \cell_outs[16] ;
 wire \cell_outs[170] ;
 wire \cell_outs[171] ;
 wire \cell_outs[172] ;
 wire \cell_outs[173] ;
 wire \cell_outs[174] ;
 wire \cell_outs[175] ;
 wire \cell_outs[176] ;
 wire \cell_outs[177] ;
 wire \cell_outs[178] ;
 wire \cell_outs[179] ;
 wire \cell_outs[17] ;
 wire \cell_outs[180] ;
 wire \cell_outs[181] ;
 wire \cell_outs[182] ;
 wire \cell_outs[183] ;
 wire \cell_outs[184] ;
 wire \cell_outs[185] ;
 wire \cell_outs[186] ;
 wire \cell_outs[187] ;
 wire \cell_outs[188] ;
 wire \cell_outs[189] ;
 wire \cell_outs[18] ;
 wire \cell_outs[190] ;
 wire \cell_outs[191] ;
 wire \cell_outs[192] ;
 wire \cell_outs[193] ;
 wire \cell_outs[194] ;
 wire \cell_outs[195] ;
 wire \cell_outs[196] ;
 wire \cell_outs[197] ;
 wire \cell_outs[198] ;
 wire \cell_outs[199] ;
 wire \cell_outs[19] ;
 wire \cell_outs[1] ;
 wire \cell_outs[200] ;
 wire \cell_outs[201] ;
 wire \cell_outs[202] ;
 wire \cell_outs[203] ;
 wire \cell_outs[204] ;
 wire \cell_outs[205] ;
 wire \cell_outs[206] ;
 wire \cell_outs[207] ;
 wire \cell_outs[208] ;
 wire \cell_outs[209] ;
 wire \cell_outs[20] ;
 wire \cell_outs[210] ;
 wire \cell_outs[211] ;
 wire \cell_outs[212] ;
 wire \cell_outs[213] ;
 wire \cell_outs[214] ;
 wire \cell_outs[215] ;
 wire \cell_outs[216] ;
 wire \cell_outs[217] ;
 wire \cell_outs[218] ;
 wire \cell_outs[219] ;
 wire \cell_outs[21] ;
 wire \cell_outs[220] ;
 wire \cell_outs[221] ;
 wire \cell_outs[222] ;
 wire \cell_outs[223] ;
 wire \cell_outs[224] ;
 wire \cell_outs[225] ;
 wire \cell_outs[226] ;
 wire \cell_outs[227] ;
 wire \cell_outs[228] ;
 wire \cell_outs[229] ;
 wire \cell_outs[22] ;
 wire \cell_outs[230] ;
 wire \cell_outs[231] ;
 wire \cell_outs[232] ;
 wire \cell_outs[233] ;
 wire \cell_outs[234] ;
 wire \cell_outs[235] ;
 wire \cell_outs[236] ;
 wire \cell_outs[237] ;
 wire \cell_outs[238] ;
 wire \cell_outs[239] ;
 wire \cell_outs[23] ;
 wire \cell_outs[240] ;
 wire \cell_outs[241] ;
 wire \cell_outs[242] ;
 wire \cell_outs[243] ;
 wire \cell_outs[244] ;
 wire \cell_outs[245] ;
 wire \cell_outs[246] ;
 wire \cell_outs[247] ;
 wire \cell_outs[248] ;
 wire \cell_outs[249] ;
 wire \cell_outs[24] ;
 wire \cell_outs[250] ;
 wire \cell_outs[251] ;
 wire \cell_outs[252] ;
 wire \cell_outs[253] ;
 wire \cell_outs[254] ;
 wire \cell_outs[255] ;
 wire \cell_outs[25] ;
 wire \cell_outs[26] ;
 wire \cell_outs[27] ;
 wire \cell_outs[28] ;
 wire \cell_outs[29] ;
 wire \cell_outs[2] ;
 wire \cell_outs[30] ;
 wire \cell_outs[31] ;
 wire \cell_outs[32] ;
 wire \cell_outs[33] ;
 wire \cell_outs[34] ;
 wire \cell_outs[35] ;
 wire \cell_outs[36] ;
 wire \cell_outs[37] ;
 wire \cell_outs[38] ;
 wire \cell_outs[39] ;
 wire \cell_outs[3] ;
 wire \cell_outs[40] ;
 wire \cell_outs[41] ;
 wire \cell_outs[42] ;
 wire \cell_outs[43] ;
 wire \cell_outs[44] ;
 wire \cell_outs[45] ;
 wire \cell_outs[46] ;
 wire \cell_outs[47] ;
 wire \cell_outs[48] ;
 wire \cell_outs[49] ;
 wire \cell_outs[4] ;
 wire \cell_outs[50] ;
 wire \cell_outs[51] ;
 wire \cell_outs[52] ;
 wire \cell_outs[53] ;
 wire \cell_outs[54] ;
 wire \cell_outs[55] ;
 wire \cell_outs[56] ;
 wire \cell_outs[57] ;
 wire \cell_outs[58] ;
 wire \cell_outs[59] ;
 wire \cell_outs[5] ;
 wire \cell_outs[60] ;
 wire \cell_outs[61] ;
 wire \cell_outs[62] ;
 wire \cell_outs[63] ;
 wire \cell_outs[64] ;
 wire \cell_outs[65] ;
 wire \cell_outs[66] ;
 wire \cell_outs[67] ;
 wire \cell_outs[68] ;
 wire \cell_outs[69] ;
 wire \cell_outs[6] ;
 wire \cell_outs[70] ;
 wire \cell_outs[71] ;
 wire \cell_outs[72] ;
 wire \cell_outs[73] ;
 wire \cell_outs[74] ;
 wire \cell_outs[75] ;
 wire \cell_outs[76] ;
 wire \cell_outs[77] ;
 wire \cell_outs[78] ;
 wire \cell_outs[79] ;
 wire \cell_outs[7] ;
 wire \cell_outs[80] ;
 wire \cell_outs[81] ;
 wire \cell_outs[82] ;
 wire \cell_outs[83] ;
 wire \cell_outs[84] ;
 wire \cell_outs[85] ;
 wire \cell_outs[86] ;
 wire \cell_outs[87] ;
 wire \cell_outs[88] ;
 wire \cell_outs[89] ;
 wire \cell_outs[8] ;
 wire \cell_outs[90] ;
 wire \cell_outs[91] ;
 wire \cell_outs[92] ;
 wire \cell_outs[93] ;
 wire \cell_outs[94] ;
 wire \cell_outs[95] ;
 wire \cell_outs[96] ;
 wire \cell_outs[97] ;
 wire \cell_outs[98] ;
 wire \cell_outs[99] ;
 wire \cell_outs[9] ;
 wire \state[0] ;
 wire \state[100] ;
 wire \state[101] ;
 wire \state[102] ;
 wire \state[103] ;
 wire \state[104] ;
 wire \state[105] ;
 wire \state[106] ;
 wire \state[107] ;
 wire \state[108] ;
 wire \state[109] ;
 wire \state[10] ;
 wire \state[110] ;
 wire \state[111] ;
 wire \state[112] ;
 wire \state[113] ;
 wire \state[114] ;
 wire \state[115] ;
 wire \state[116] ;
 wire \state[117] ;
 wire \state[118] ;
 wire \state[119] ;
 wire \state[11] ;
 wire \state[120] ;
 wire \state[121] ;
 wire \state[122] ;
 wire \state[123] ;
 wire \state[124] ;
 wire \state[125] ;
 wire \state[126] ;
 wire \state[127] ;
 wire \state[128] ;
 wire \state[129] ;
 wire \state[12] ;
 wire \state[130] ;
 wire \state[131] ;
 wire \state[132] ;
 wire \state[133] ;
 wire \state[134] ;
 wire \state[135] ;
 wire \state[136] ;
 wire \state[137] ;
 wire \state[138] ;
 wire \state[139] ;
 wire \state[13] ;
 wire \state[140] ;
 wire \state[141] ;
 wire \state[142] ;
 wire \state[143] ;
 wire \state[144] ;
 wire \state[145] ;
 wire \state[146] ;
 wire \state[147] ;
 wire \state[148] ;
 wire \state[149] ;
 wire \state[14] ;
 wire \state[150] ;
 wire \state[151] ;
 wire \state[152] ;
 wire \state[153] ;
 wire \state[154] ;
 wire \state[155] ;
 wire \state[156] ;
 wire \state[157] ;
 wire \state[158] ;
 wire \state[159] ;
 wire \state[15] ;
 wire \state[160] ;
 wire \state[161] ;
 wire \state[162] ;
 wire \state[163] ;
 wire \state[164] ;
 wire \state[165] ;
 wire \state[166] ;
 wire \state[167] ;
 wire \state[168] ;
 wire \state[169] ;
 wire \state[16] ;
 wire \state[170] ;
 wire \state[171] ;
 wire \state[172] ;
 wire \state[173] ;
 wire \state[174] ;
 wire \state[175] ;
 wire \state[176] ;
 wire \state[177] ;
 wire \state[178] ;
 wire \state[179] ;
 wire \state[17] ;
 wire \state[180] ;
 wire \state[181] ;
 wire \state[182] ;
 wire \state[183] ;
 wire \state[184] ;
 wire \state[185] ;
 wire \state[186] ;
 wire \state[187] ;
 wire \state[188] ;
 wire \state[189] ;
 wire \state[18] ;
 wire \state[190] ;
 wire \state[191] ;
 wire \state[192] ;
 wire \state[193] ;
 wire \state[194] ;
 wire \state[195] ;
 wire \state[196] ;
 wire \state[197] ;
 wire \state[198] ;
 wire \state[199] ;
 wire \state[19] ;
 wire \state[1] ;
 wire \state[200] ;
 wire \state[201] ;
 wire \state[202] ;
 wire \state[203] ;
 wire \state[204] ;
 wire \state[205] ;
 wire \state[206] ;
 wire \state[207] ;
 wire \state[208] ;
 wire \state[209] ;
 wire \state[20] ;
 wire \state[210] ;
 wire \state[211] ;
 wire \state[212] ;
 wire \state[213] ;
 wire \state[214] ;
 wire \state[215] ;
 wire \state[216] ;
 wire \state[217] ;
 wire \state[218] ;
 wire \state[219] ;
 wire \state[21] ;
 wire \state[220] ;
 wire \state[221] ;
 wire \state[222] ;
 wire \state[223] ;
 wire \state[224] ;
 wire \state[225] ;
 wire \state[226] ;
 wire \state[227] ;
 wire \state[228] ;
 wire \state[229] ;
 wire \state[22] ;
 wire \state[230] ;
 wire \state[231] ;
 wire \state[232] ;
 wire \state[233] ;
 wire \state[234] ;
 wire \state[235] ;
 wire \state[236] ;
 wire \state[237] ;
 wire \state[238] ;
 wire \state[239] ;
 wire \state[23] ;
 wire \state[240] ;
 wire \state[241] ;
 wire \state[242] ;
 wire \state[243] ;
 wire \state[244] ;
 wire \state[245] ;
 wire \state[246] ;
 wire \state[247] ;
 wire \state[248] ;
 wire \state[249] ;
 wire \state[24] ;
 wire \state[250] ;
 wire \state[251] ;
 wire \state[252] ;
 wire \state[253] ;
 wire \state[254] ;
 wire \state[255] ;
 wire \state[25] ;
 wire \state[26] ;
 wire \state[27] ;
 wire \state[28] ;
 wire \state[29] ;
 wire \state[2] ;
 wire \state[30] ;
 wire \state[31] ;
 wire \state[32] ;
 wire \state[33] ;
 wire \state[34] ;
 wire \state[35] ;
 wire \state[36] ;
 wire \state[37] ;
 wire \state[38] ;
 wire \state[39] ;
 wire \state[3] ;
 wire \state[40] ;
 wire \state[41] ;
 wire \state[42] ;
 wire \state[43] ;
 wire \state[44] ;
 wire \state[45] ;
 wire \state[46] ;
 wire \state[47] ;
 wire \state[48] ;
 wire \state[49] ;
 wire \state[4] ;
 wire \state[50] ;
 wire \state[51] ;
 wire \state[52] ;
 wire \state[53] ;
 wire \state[54] ;
 wire \state[55] ;
 wire \state[56] ;
 wire \state[57] ;
 wire \state[58] ;
 wire \state[59] ;
 wire \state[5] ;
 wire \state[60] ;
 wire \state[61] ;
 wire \state[62] ;
 wire \state[63] ;
 wire \state[64] ;
 wire \state[65] ;
 wire \state[66] ;
 wire \state[67] ;
 wire \state[68] ;
 wire \state[69] ;
 wire \state[6] ;
 wire \state[70] ;
 wire \state[71] ;
 wire \state[72] ;
 wire \state[73] ;
 wire \state[74] ;
 wire \state[75] ;
 wire \state[76] ;
 wire \state[77] ;
 wire \state[78] ;
 wire \state[79] ;
 wire \state[7] ;
 wire \state[80] ;
 wire \state[81] ;
 wire \state[82] ;
 wire \state[83] ;
 wire \state[84] ;
 wire \state[85] ;
 wire \state[86] ;
 wire \state[87] ;
 wire \state[88] ;
 wire \state[89] ;
 wire \state[8] ;
 wire \state[90] ;
 wire \state[91] ;
 wire \state[92] ;
 wire \state[93] ;
 wire \state[94] ;
 wire \state[95] ;
 wire \state[96] ;
 wire \state[97] ;
 wire \state[98] ;
 wire \state[99] ;
 wire \state[9] ;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net327;

 sky130_fd_sc_hd__or3_2 _34_ (.A(net116),
    .B(net118),
    .C(net120),
    .X(_16_));
 sky130_fd_sc_hd__nor3b_2 _35_ (.A(_16_),
    .B(net21),
    .C_N(net17),
    .Y(_01_));
 sky130_fd_sc_hd__and2b_2 _36_ (.A_N(net21),
    .B(net17),
    .X(_17_));
 sky130_fd_sc_hd__and4bb_2 _37_ (.A_N(net116),
    .B_N(net118),
    .C(net120),
    .D(_17_),
    .X(_18_));
 sky130_fd_sc_hd__buf_12 _38_ (.A(_18_),
    .X(_11_));
 sky130_fd_sc_hd__and4bb_2 _39_ (.A_N(net116),
    .B_N(net120),
    .C(_17_),
    .D(net118),
    .X(_19_));
 sky130_fd_sc_hd__buf_12 _40_ (.A(_19_),
    .X(_00_));
 sky130_fd_sc_hd__and4b_1 _41_ (.A_N(net116),
    .B(net118),
    .C(net120),
    .D(_17_),
    .X(_20_));
 sky130_fd_sc_hd__buf_12 _42_ (.A(_20_),
    .X(_02_));
 sky130_fd_sc_hd__and4bb_1 _43_ (.A_N(net118),
    .B_N(net120),
    .C(_17_),
    .D(net116),
    .X(_21_));
 sky130_fd_sc_hd__buf_12 _44_ (.A(_21_),
    .X(_03_));
 sky130_fd_sc_hd__and4b_1 _45_ (.A_N(net118),
    .B(net120),
    .C(_17_),
    .D(net116),
    .X(_22_));
 sky130_fd_sc_hd__buf_12 _46_ (.A(_22_),
    .X(_04_));
 sky130_fd_sc_hd__and4b_1 _47_ (.A_N(net120),
    .B(_17_),
    .C(net116),
    .D(net118),
    .X(_23_));
 sky130_fd_sc_hd__buf_12 _48_ (.A(_23_),
    .X(_05_));
 sky130_fd_sc_hd__and4_1 _49_ (.A(net116),
    .B(net118),
    .C(net120),
    .D(_17_),
    .X(_24_));
 sky130_fd_sc_hd__buf_12 _50_ (.A(_24_),
    .X(_06_));
 sky130_fd_sc_hd__and2_4 _51_ (.A(net21),
    .B(net17),
    .X(_25_));
 sky130_fd_sc_hd__and2b_1 _52_ (.A_N(_16_),
    .B(_25_),
    .X(_26_));
 sky130_fd_sc_hd__buf_12 _53_ (.A(_26_),
    .X(_07_));
 sky130_fd_sc_hd__and4bb_1 _54_ (.A_N(net116),
    .B_N(net118),
    .C(net120),
    .D(_25_),
    .X(_27_));
 sky130_fd_sc_hd__buf_12 _55_ (.A(_27_),
    .X(_08_));
 sky130_fd_sc_hd__and4bb_1 _56_ (.A_N(net116),
    .B_N(net120),
    .C(_25_),
    .D(net118),
    .X(_28_));
 sky130_fd_sc_hd__buf_12 _57_ (.A(_28_),
    .X(_09_));
 sky130_fd_sc_hd__and4b_1 _58_ (.A_N(net117),
    .B(net119),
    .C(net121),
    .D(_25_),
    .X(_29_));
 sky130_fd_sc_hd__buf_12 _59_ (.A(_29_),
    .X(_10_));
 sky130_fd_sc_hd__and4bb_1 _60_ (.A_N(net119),
    .B_N(net121),
    .C(_25_),
    .D(net117),
    .X(_30_));
 sky130_fd_sc_hd__buf_12 _61_ (.A(_30_),
    .X(_12_));
 sky130_fd_sc_hd__and4b_1 _62_ (.A_N(net119),
    .B(net121),
    .C(_25_),
    .D(net117),
    .X(_31_));
 sky130_fd_sc_hd__buf_12 _63_ (.A(_31_),
    .X(_13_));
 sky130_fd_sc_hd__and4b_1 _64_ (.A_N(net121),
    .B(_25_),
    .C(net117),
    .D(net119),
    .X(_32_));
 sky130_fd_sc_hd__buf_12 _65_ (.A(_32_),
    .X(_14_));
 sky130_fd_sc_hd__and4_2 _66_ (.A(net117),
    .B(net119),
    .C(net121),
    .D(_25_),
    .X(_33_));
 sky130_fd_sc_hd__buf_12 _67_ (.A(_33_),
    .X(_15_));
 sky130_fd_sc_hd__clkbuf_2 _68_ (.A(\cell_outs[0] ),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 _69_ (.A(\cell_outs[1] ),
    .X(net33));
 sky130_fd_sc_hd__buf_1 _70_ (.A(\cell_outs[2] ),
    .X(net34));
 sky130_fd_sc_hd__buf_1 _71_ (.A(\cell_outs[3] ),
    .X(net35));
 sky130_fd_sc_hd__buf_8 _72_ (.A(\cell_outs[4] ),
    .X(net36));
 sky130_fd_sc_hd__buf_1 _73_ (.A(\cell_outs[5] ),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_8 _74_ (.A(net49),
    .X(net38));
 sky130_fd_sc_hd__buf_12 _75_ (.A(\cell_outs[7] ),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_16 _76_ (.A(\cell_outs[8] ),
    .X(net40));
 sky130_fd_sc_hd__buf_8 _77_ (.A(\cell_outs[9] ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 _78_ (.A(\cell_outs[10] ),
    .X(net27));
 sky130_fd_sc_hd__buf_12 _79_ (.A(\cell_outs[11] ),
    .X(net28));
 sky130_fd_sc_hd__buf_6 _80_ (.A(\cell_outs[12] ),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 _81_ (.A(\cell_outs[13] ),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_16 _82_ (.A(\cell_outs[14] ),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 _83_ (.A(\cell_outs[15] ),
    .X(net32));
 life_cell arr_cell_x0_y0 (.clk(clknet_5_0__leaf_clk),
    .d(net123),
    .dl(net124),
    .dr(net125),
    .in_data(net122),
    .l(net126),
    .load_in(net42),
    .load_out(net22),
    .out_data(\cell_outs[0] ),
    .prev_out_data(\cell_outs[16] ),
    .r(\state[1] ),
    .reset(net24),
    .run(net52),
    .shift(net23),
    .state(\state[0] ),
    .u(\state[16] ),
    .ul(net127),
    .ur(\state[17] ));
 life_cell arr_cell_x0_y1 (.clk(clknet_5_0__leaf_clk),
    .d(\state[0] ),
    .dl(net128),
    .dr(\state[1] ),
    .in_data(net122),
    .l(net129),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[16] ),
    .prev_out_data(\cell_outs[32] ),
    .r(\state[17] ),
    .reset(net24),
    .run(net53),
    .shift(net23),
    .state(\state[16] ),
    .u(\state[32] ),
    .ul(net130),
    .ur(\state[33] ));
 life_cell arr_cell_x0_y10 (.clk(clknet_5_17__leaf_clk),
    .d(\state[144] ),
    .dl(net131),
    .dr(\state[145] ),
    .in_data(net122),
    .l(net132),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[160] ),
    .prev_out_data(\cell_outs[176] ),
    .r(\state[161] ),
    .reset(net24),
    .run(net63),
    .shift(net23),
    .state(\state[160] ),
    .u(\state[176] ),
    .ul(net133),
    .ur(\state[177] ));
 life_cell arr_cell_x0_y11 (.clk(clknet_5_17__leaf_clk),
    .d(\state[160] ),
    .dl(net134),
    .dr(\state[161] ),
    .in_data(net122),
    .l(net135),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[176] ),
    .prev_out_data(\cell_outs[192] ),
    .r(\state[177] ),
    .reset(net24),
    .run(net62),
    .shift(net23),
    .state(\state[176] ),
    .u(\state[192] ),
    .ul(net136),
    .ur(\state[193] ));
 life_cell arr_cell_x0_y12 (.clk(clknet_5_20__leaf_clk),
    .d(\state[176] ),
    .dl(net137),
    .dr(\state[177] ),
    .in_data(net122),
    .l(net138),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[192] ),
    .prev_out_data(\cell_outs[208] ),
    .r(\state[193] ),
    .reset(net24),
    .run(net61),
    .shift(net23),
    .state(\state[192] ),
    .u(\state[208] ),
    .ul(net139),
    .ur(\state[209] ));
 life_cell arr_cell_x0_y13 (.clk(clknet_5_20__leaf_clk),
    .d(\state[192] ),
    .dl(net140),
    .dr(\state[193] ),
    .in_data(net122),
    .l(net141),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[208] ),
    .prev_out_data(\cell_outs[224] ),
    .r(\state[209] ),
    .reset(net24),
    .run(net60),
    .shift(net23),
    .state(\state[208] ),
    .u(\state[224] ),
    .ul(net142),
    .ur(\state[225] ));
 life_cell arr_cell_x0_y14 (.clk(clknet_5_21__leaf_clk),
    .d(\state[208] ),
    .dl(net143),
    .dr(\state[209] ),
    .in_data(net122),
    .l(net144),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[224] ),
    .prev_out_data(\cell_outs[240] ),
    .r(\state[225] ),
    .reset(net24),
    .run(net59),
    .shift(net23),
    .state(\state[224] ),
    .u(\state[240] ),
    .ul(net145),
    .ur(\state[241] ));
 life_cell arr_cell_x0_y15 (.clk(clknet_5_21__leaf_clk),
    .d(\state[224] ),
    .dl(net146),
    .dr(\state[225] ),
    .in_data(net122),
    .l(net147),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[240] ),
    .prev_out_data(net148),
    .r(\state[241] ),
    .reset(net24),
    .run(net58),
    .shift(net23),
    .state(\state[240] ),
    .u(net149),
    .ul(net150),
    .ur(net151));
 life_cell arr_cell_x0_y2 (.clk(clknet_5_1__leaf_clk),
    .d(\state[16] ),
    .dl(net152),
    .dr(\state[17] ),
    .in_data(net122),
    .l(net153),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[32] ),
    .prev_out_data(\cell_outs[48] ),
    .r(\state[33] ),
    .reset(net24),
    .run(net54),
    .shift(net23),
    .state(\state[32] ),
    .u(\state[48] ),
    .ul(net154),
    .ur(\state[49] ));
 life_cell arr_cell_x0_y3 (.clk(clknet_5_1__leaf_clk),
    .d(\state[32] ),
    .dl(net155),
    .dr(\state[33] ),
    .in_data(net122),
    .l(net156),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[48] ),
    .prev_out_data(\cell_outs[64] ),
    .r(\state[49] ),
    .reset(net24),
    .run(net55),
    .shift(net23),
    .state(\state[48] ),
    .u(\state[64] ),
    .ul(net157),
    .ur(\state[65] ));
 life_cell arr_cell_x0_y4 (.clk(clknet_5_4__leaf_clk),
    .d(\state[48] ),
    .dl(net158),
    .dr(\state[49] ),
    .in_data(net122),
    .l(net159),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[64] ),
    .prev_out_data(\cell_outs[80] ),
    .r(\state[65] ),
    .reset(net24),
    .run(net56),
    .shift(net23),
    .state(\state[64] ),
    .u(\state[80] ),
    .ul(net160),
    .ur(\state[81] ));
 life_cell arr_cell_x0_y5 (.clk(clknet_5_4__leaf_clk),
    .d(\state[64] ),
    .dl(net161),
    .dr(\state[65] ),
    .in_data(net122),
    .l(net162),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[80] ),
    .prev_out_data(\cell_outs[96] ),
    .r(\state[81] ),
    .reset(net24),
    .run(net57),
    .shift(net23),
    .state(\state[80] ),
    .u(\state[96] ),
    .ul(net163),
    .ur(\state[97] ));
 life_cell arr_cell_x0_y6 (.clk(clknet_5_5__leaf_clk),
    .d(\state[80] ),
    .dl(net164),
    .dr(\state[81] ),
    .in_data(net122),
    .l(net165),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[96] ),
    .prev_out_data(\cell_outs[112] ),
    .r(\state[97] ),
    .reset(net24),
    .run(net66),
    .shift(net23),
    .state(\state[96] ),
    .u(\state[112] ),
    .ul(net166),
    .ur(\state[113] ));
 life_cell arr_cell_x0_y7 (.clk(clknet_5_5__leaf_clk),
    .d(\state[96] ),
    .dl(net167),
    .dr(\state[97] ),
    .in_data(net122),
    .l(net168),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[112] ),
    .prev_out_data(\cell_outs[128] ),
    .r(\state[113] ),
    .reset(net24),
    .run(net25),
    .shift(net23),
    .state(\state[112] ),
    .u(\state[128] ),
    .ul(net169),
    .ur(\state[129] ));
 life_cell arr_cell_x0_y8 (.clk(clknet_5_16__leaf_clk),
    .d(\state[112] ),
    .dl(net170),
    .dr(\state[113] ),
    .in_data(net122),
    .l(net171),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[128] ),
    .prev_out_data(\cell_outs[144] ),
    .r(\state[129] ),
    .reset(net24),
    .run(net65),
    .shift(net23),
    .state(\state[128] ),
    .u(\state[144] ),
    .ul(net172),
    .ur(\state[145] ));
 life_cell arr_cell_x0_y9 (.clk(clknet_5_16__leaf_clk),
    .d(\state[128] ),
    .dl(net173),
    .dr(\state[129] ),
    .in_data(net122),
    .l(net174),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[144] ),
    .prev_out_data(\cell_outs[160] ),
    .r(\state[145] ),
    .reset(net24),
    .run(net64),
    .shift(net23),
    .state(\state[144] ),
    .u(\state[160] ),
    .ul(net175),
    .ur(\state[161] ));
 life_cell arr_cell_x10_y0 (.clk(clknet_5_8__leaf_clk),
    .d(net176),
    .dl(net177),
    .dr(net178),
    .in_data(net2),
    .l(\state[9] ),
    .load_in(net45),
    .load_out(net22),
    .out_data(\cell_outs[10] ),
    .prev_out_data(\cell_outs[26] ),
    .r(\state[11] ),
    .reset(net72),
    .run(net52),
    .shift(net87),
    .state(\state[10] ),
    .u(\state[26] ),
    .ul(\state[25] ),
    .ur(\state[27] ));
 life_cell arr_cell_x10_y1 (.clk(clknet_5_8__leaf_clk),
    .d(\state[10] ),
    .dl(\state[9] ),
    .dr(\state[11] ),
    .in_data(net2),
    .l(\state[25] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[26] ),
    .prev_out_data(\cell_outs[42] ),
    .r(\state[27] ),
    .reset(net72),
    .run(net53),
    .shift(net87),
    .state(\state[26] ),
    .u(\state[42] ),
    .ul(\state[41] ),
    .ur(\state[43] ));
 life_cell arr_cell_x10_y10 (.clk(clknet_5_25__leaf_clk),
    .d(\state[154] ),
    .dl(\state[153] ),
    .dr(\state[155] ),
    .in_data(net2),
    .l(\state[169] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[170] ),
    .prev_out_data(\cell_outs[186] ),
    .r(\state[171] ),
    .reset(net72),
    .run(net63),
    .shift(net87),
    .state(\state[170] ),
    .u(\state[186] ),
    .ul(\state[185] ),
    .ur(\state[187] ));
 life_cell arr_cell_x10_y11 (.clk(clknet_5_25__leaf_clk),
    .d(\state[170] ),
    .dl(\state[169] ),
    .dr(\state[171] ),
    .in_data(net2),
    .l(\state[185] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[186] ),
    .prev_out_data(\cell_outs[202] ),
    .r(\state[187] ),
    .reset(net72),
    .run(net62),
    .shift(net87),
    .state(\state[186] ),
    .u(\state[202] ),
    .ul(\state[201] ),
    .ur(\state[203] ));
 life_cell arr_cell_x10_y12 (.clk(clknet_5_28__leaf_clk),
    .d(\state[186] ),
    .dl(\state[185] ),
    .dr(\state[187] ),
    .in_data(net2),
    .l(\state[201] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[202] ),
    .prev_out_data(\cell_outs[218] ),
    .r(\state[203] ),
    .reset(net72),
    .run(net61),
    .shift(net87),
    .state(\state[202] ),
    .u(\state[218] ),
    .ul(\state[217] ),
    .ur(\state[219] ));
 life_cell arr_cell_x10_y13 (.clk(clknet_5_28__leaf_clk),
    .d(\state[202] ),
    .dl(\state[201] ),
    .dr(\state[203] ),
    .in_data(net2),
    .l(\state[217] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[218] ),
    .prev_out_data(\cell_outs[234] ),
    .r(\state[219] ),
    .reset(net72),
    .run(net60),
    .shift(net87),
    .state(\state[218] ),
    .u(\state[234] ),
    .ul(\state[233] ),
    .ur(\state[235] ));
 life_cell arr_cell_x10_y14 (.clk(clknet_5_29__leaf_clk),
    .d(\state[218] ),
    .dl(\state[217] ),
    .dr(\state[219] ),
    .in_data(net2),
    .l(\state[233] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[234] ),
    .prev_out_data(\cell_outs[250] ),
    .r(\state[235] ),
    .reset(net72),
    .run(net59),
    .shift(net87),
    .state(\state[234] ),
    .u(\state[250] ),
    .ul(\state[249] ),
    .ur(\state[251] ));
 life_cell arr_cell_x10_y15 (.clk(clknet_5_29__leaf_clk),
    .d(\state[234] ),
    .dl(\state[233] ),
    .dr(\state[235] ),
    .in_data(net2),
    .l(\state[249] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[250] ),
    .prev_out_data(net179),
    .r(\state[251] ),
    .reset(net72),
    .run(net58),
    .shift(net87),
    .state(\state[250] ),
    .u(net180),
    .ul(net181),
    .ur(net182));
 life_cell arr_cell_x10_y2 (.clk(clknet_5_9__leaf_clk),
    .d(\state[26] ),
    .dl(\state[25] ),
    .dr(\state[27] ),
    .in_data(net2),
    .l(\state[41] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[42] ),
    .prev_out_data(\cell_outs[58] ),
    .r(\state[43] ),
    .reset(net72),
    .run(net54),
    .shift(net87),
    .state(\state[42] ),
    .u(\state[58] ),
    .ul(\state[57] ),
    .ur(\state[59] ));
 life_cell arr_cell_x10_y3 (.clk(clknet_5_9__leaf_clk),
    .d(\state[42] ),
    .dl(\state[41] ),
    .dr(\state[43] ),
    .in_data(net2),
    .l(\state[57] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[58] ),
    .prev_out_data(\cell_outs[74] ),
    .r(\state[59] ),
    .reset(net72),
    .run(net55),
    .shift(net87),
    .state(\state[58] ),
    .u(\state[74] ),
    .ul(\state[73] ),
    .ur(\state[75] ));
 life_cell arr_cell_x10_y4 (.clk(clknet_5_12__leaf_clk),
    .d(\state[58] ),
    .dl(\state[57] ),
    .dr(\state[59] ),
    .in_data(net2),
    .l(\state[73] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[74] ),
    .prev_out_data(\cell_outs[90] ),
    .r(\state[75] ),
    .reset(net72),
    .run(net56),
    .shift(net87),
    .state(\state[74] ),
    .u(\state[90] ),
    .ul(\state[89] ),
    .ur(\state[91] ));
 life_cell arr_cell_x10_y5 (.clk(clknet_5_12__leaf_clk),
    .d(\state[74] ),
    .dl(\state[73] ),
    .dr(\state[75] ),
    .in_data(net2),
    .l(\state[89] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[90] ),
    .prev_out_data(\cell_outs[106] ),
    .r(\state[91] ),
    .reset(net72),
    .run(net57),
    .shift(net87),
    .state(\state[90] ),
    .u(\state[106] ),
    .ul(\state[105] ),
    .ur(\state[107] ));
 life_cell arr_cell_x10_y6 (.clk(clknet_5_13__leaf_clk),
    .d(\state[90] ),
    .dl(\state[89] ),
    .dr(\state[91] ),
    .in_data(net2),
    .l(\state[105] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[106] ),
    .prev_out_data(\cell_outs[122] ),
    .r(\state[107] ),
    .reset(net72),
    .run(net66),
    .shift(net87),
    .state(\state[106] ),
    .u(\state[122] ),
    .ul(\state[121] ),
    .ur(\state[123] ));
 life_cell arr_cell_x10_y7 (.clk(clknet_5_13__leaf_clk),
    .d(\state[106] ),
    .dl(\state[105] ),
    .dr(\state[107] ),
    .in_data(net2),
    .l(\state[121] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[122] ),
    .prev_out_data(\cell_outs[138] ),
    .r(\state[123] ),
    .reset(net72),
    .run(net25),
    .shift(net87),
    .state(\state[122] ),
    .u(\state[138] ),
    .ul(\state[137] ),
    .ur(\state[139] ));
 life_cell arr_cell_x10_y8 (.clk(clknet_5_24__leaf_clk),
    .d(\state[122] ),
    .dl(\state[121] ),
    .dr(\state[123] ),
    .in_data(net2),
    .l(\state[137] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[138] ),
    .prev_out_data(\cell_outs[154] ),
    .r(\state[139] ),
    .reset(net72),
    .run(net65),
    .shift(net87),
    .state(\state[138] ),
    .u(\state[154] ),
    .ul(\state[153] ),
    .ur(\state[155] ));
 life_cell arr_cell_x10_y9 (.clk(clknet_5_24__leaf_clk),
    .d(\state[138] ),
    .dl(\state[137] ),
    .dr(\state[139] ),
    .in_data(net2),
    .l(\state[153] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[154] ),
    .prev_out_data(\cell_outs[170] ),
    .r(\state[155] ),
    .reset(net72),
    .run(net64),
    .shift(net87),
    .state(\state[154] ),
    .u(\state[170] ),
    .ul(\state[169] ),
    .ur(\state[171] ));
 life_cell arr_cell_x11_y0 (.clk(clknet_5_8__leaf_clk),
    .d(net183),
    .dl(net184),
    .dr(net185),
    .in_data(net3),
    .l(\state[10] ),
    .load_in(net44),
    .load_out(net115),
    .out_data(\cell_outs[11] ),
    .prev_out_data(\cell_outs[27] ),
    .r(\state[12] ),
    .reset(net71),
    .run(net52),
    .shift(net86),
    .state(\state[11] ),
    .u(\state[27] ),
    .ul(\state[26] ),
    .ur(\state[28] ));
 life_cell arr_cell_x11_y1 (.clk(clknet_5_8__leaf_clk),
    .d(\state[11] ),
    .dl(\state[10] ),
    .dr(\state[12] ),
    .in_data(net3),
    .l(\state[26] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[27] ),
    .prev_out_data(\cell_outs[43] ),
    .r(\state[28] ),
    .reset(net71),
    .run(net53),
    .shift(net86),
    .state(\state[27] ),
    .u(\state[43] ),
    .ul(\state[42] ),
    .ur(\state[44] ));
 life_cell arr_cell_x11_y10 (.clk(clknet_5_25__leaf_clk),
    .d(\state[155] ),
    .dl(\state[154] ),
    .dr(\state[156] ),
    .in_data(net3),
    .l(\state[170] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[171] ),
    .prev_out_data(\cell_outs[187] ),
    .r(\state[172] ),
    .reset(net71),
    .run(net63),
    .shift(net86),
    .state(\state[171] ),
    .u(\state[187] ),
    .ul(\state[186] ),
    .ur(\state[188] ));
 life_cell arr_cell_x11_y11 (.clk(clknet_5_25__leaf_clk),
    .d(\state[171] ),
    .dl(\state[170] ),
    .dr(\state[172] ),
    .in_data(net3),
    .l(\state[186] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[187] ),
    .prev_out_data(\cell_outs[203] ),
    .r(\state[188] ),
    .reset(net71),
    .run(net62),
    .shift(net86),
    .state(\state[187] ),
    .u(\state[203] ),
    .ul(\state[202] ),
    .ur(\state[204] ));
 life_cell arr_cell_x11_y12 (.clk(clknet_5_28__leaf_clk),
    .d(\state[187] ),
    .dl(\state[186] ),
    .dr(\state[188] ),
    .in_data(net3),
    .l(\state[202] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[203] ),
    .prev_out_data(\cell_outs[219] ),
    .r(\state[204] ),
    .reset(net71),
    .run(net61),
    .shift(net86),
    .state(\state[203] ),
    .u(\state[219] ),
    .ul(\state[218] ),
    .ur(\state[220] ));
 life_cell arr_cell_x11_y13 (.clk(clknet_5_28__leaf_clk),
    .d(\state[203] ),
    .dl(\state[202] ),
    .dr(\state[204] ),
    .in_data(net3),
    .l(\state[218] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[219] ),
    .prev_out_data(\cell_outs[235] ),
    .r(\state[220] ),
    .reset(net71),
    .run(net60),
    .shift(net86),
    .state(\state[219] ),
    .u(\state[235] ),
    .ul(\state[234] ),
    .ur(\state[236] ));
 life_cell arr_cell_x11_y14 (.clk(clknet_5_29__leaf_clk),
    .d(\state[219] ),
    .dl(\state[218] ),
    .dr(\state[220] ),
    .in_data(net3),
    .l(\state[234] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[235] ),
    .prev_out_data(\cell_outs[251] ),
    .r(\state[236] ),
    .reset(net71),
    .run(net59),
    .shift(net86),
    .state(\state[235] ),
    .u(\state[251] ),
    .ul(\state[250] ),
    .ur(\state[252] ));
 life_cell arr_cell_x11_y15 (.clk(clknet_5_29__leaf_clk),
    .d(\state[235] ),
    .dl(\state[234] ),
    .dr(\state[236] ),
    .in_data(net3),
    .l(\state[250] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[251] ),
    .prev_out_data(net186),
    .r(\state[252] ),
    .reset(net71),
    .run(net58),
    .shift(net86),
    .state(\state[251] ),
    .u(net187),
    .ul(net188),
    .ur(net189));
 life_cell arr_cell_x11_y2 (.clk(clknet_5_9__leaf_clk),
    .d(\state[27] ),
    .dl(\state[26] ),
    .dr(\state[28] ),
    .in_data(net3),
    .l(\state[42] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[43] ),
    .prev_out_data(\cell_outs[59] ),
    .r(\state[44] ),
    .reset(net71),
    .run(net54),
    .shift(net86),
    .state(\state[43] ),
    .u(\state[59] ),
    .ul(\state[58] ),
    .ur(\state[60] ));
 life_cell arr_cell_x11_y3 (.clk(clknet_5_9__leaf_clk),
    .d(\state[43] ),
    .dl(\state[42] ),
    .dr(\state[44] ),
    .in_data(net3),
    .l(\state[58] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[59] ),
    .prev_out_data(\cell_outs[75] ),
    .r(\state[60] ),
    .reset(net71),
    .run(net55),
    .shift(net86),
    .state(\state[59] ),
    .u(\state[75] ),
    .ul(\state[74] ),
    .ur(\state[76] ));
 life_cell arr_cell_x11_y4 (.clk(clknet_5_12__leaf_clk),
    .d(\state[59] ),
    .dl(\state[58] ),
    .dr(\state[60] ),
    .in_data(net3),
    .l(\state[74] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[75] ),
    .prev_out_data(\cell_outs[91] ),
    .r(\state[76] ),
    .reset(net71),
    .run(net56),
    .shift(net86),
    .state(\state[75] ),
    .u(\state[91] ),
    .ul(\state[90] ),
    .ur(\state[92] ));
 life_cell arr_cell_x11_y5 (.clk(clknet_5_12__leaf_clk),
    .d(\state[75] ),
    .dl(\state[74] ),
    .dr(\state[76] ),
    .in_data(net3),
    .l(\state[90] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[91] ),
    .prev_out_data(\cell_outs[107] ),
    .r(\state[92] ),
    .reset(net71),
    .run(net57),
    .shift(net86),
    .state(\state[91] ),
    .u(\state[107] ),
    .ul(\state[106] ),
    .ur(\state[108] ));
 life_cell arr_cell_x11_y6 (.clk(clknet_5_13__leaf_clk),
    .d(\state[91] ),
    .dl(\state[90] ),
    .dr(\state[92] ),
    .in_data(net3),
    .l(\state[106] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[107] ),
    .prev_out_data(\cell_outs[123] ),
    .r(\state[108] ),
    .reset(net71),
    .run(net66),
    .shift(net86),
    .state(\state[107] ),
    .u(\state[123] ),
    .ul(\state[122] ),
    .ur(\state[124] ));
 life_cell arr_cell_x11_y7 (.clk(clknet_5_13__leaf_clk),
    .d(\state[107] ),
    .dl(\state[106] ),
    .dr(\state[108] ),
    .in_data(net3),
    .l(\state[122] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[123] ),
    .prev_out_data(\cell_outs[139] ),
    .r(\state[124] ),
    .reset(net71),
    .run(net25),
    .shift(net86),
    .state(\state[123] ),
    .u(\state[139] ),
    .ul(\state[138] ),
    .ur(\state[140] ));
 life_cell arr_cell_x11_y8 (.clk(clknet_5_24__leaf_clk),
    .d(\state[123] ),
    .dl(\state[122] ),
    .dr(\state[124] ),
    .in_data(net3),
    .l(\state[138] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[139] ),
    .prev_out_data(\cell_outs[155] ),
    .r(\state[140] ),
    .reset(net71),
    .run(net65),
    .shift(net86),
    .state(\state[139] ),
    .u(\state[155] ),
    .ul(\state[154] ),
    .ur(\state[156] ));
 life_cell arr_cell_x11_y9 (.clk(clknet_5_24__leaf_clk),
    .d(\state[139] ),
    .dl(\state[138] ),
    .dr(\state[140] ),
    .in_data(net3),
    .l(\state[154] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[155] ),
    .prev_out_data(\cell_outs[171] ),
    .r(\state[156] ),
    .reset(net71),
    .run(net64),
    .shift(net86),
    .state(\state[155] ),
    .u(\state[171] ),
    .ul(\state[170] ),
    .ur(\state[172] ));
 life_cell arr_cell_x12_y0 (.clk(clknet_5_10__leaf_clk),
    .d(net190),
    .dl(net191),
    .dr(net192),
    .in_data(net4),
    .l(\state[11] ),
    .load_in(net44),
    .load_out(net114),
    .out_data(\cell_outs[12] ),
    .prev_out_data(\cell_outs[28] ),
    .r(\state[13] ),
    .reset(net70),
    .run(net52),
    .shift(net85),
    .state(\state[12] ),
    .u(\state[28] ),
    .ul(\state[27] ),
    .ur(\state[29] ));
 life_cell arr_cell_x12_y1 (.clk(clknet_5_10__leaf_clk),
    .d(\state[12] ),
    .dl(\state[11] ),
    .dr(\state[13] ),
    .in_data(net4),
    .l(\state[27] ),
    .load_in(_11_),
    .load_out(net114),
    .out_data(\cell_outs[28] ),
    .prev_out_data(\cell_outs[44] ),
    .r(\state[29] ),
    .reset(net70),
    .run(net53),
    .shift(net85),
    .state(\state[28] ),
    .u(\state[44] ),
    .ul(\state[43] ),
    .ur(\state[45] ));
 life_cell arr_cell_x12_y10 (.clk(clknet_5_27__leaf_clk),
    .d(\state[156] ),
    .dl(\state[155] ),
    .dr(\state[157] ),
    .in_data(net4),
    .l(\state[171] ),
    .load_in(_09_),
    .load_out(net114),
    .out_data(\cell_outs[172] ),
    .prev_out_data(\cell_outs[188] ),
    .r(\state[173] ),
    .reset(net70),
    .run(net63),
    .shift(net85),
    .state(\state[172] ),
    .u(\state[188] ),
    .ul(\state[187] ),
    .ur(\state[189] ));
 life_cell arr_cell_x12_y11 (.clk(clknet_5_27__leaf_clk),
    .d(\state[172] ),
    .dl(\state[171] ),
    .dr(\state[173] ),
    .in_data(net4),
    .l(\state[187] ),
    .load_in(_10_),
    .load_out(net114),
    .out_data(\cell_outs[188] ),
    .prev_out_data(\cell_outs[204] ),
    .r(\state[189] ),
    .reset(net70),
    .run(net62),
    .shift(net85),
    .state(\state[188] ),
    .u(\state[204] ),
    .ul(\state[203] ),
    .ur(\state[205] ));
 life_cell arr_cell_x12_y12 (.clk(clknet_5_30__leaf_clk),
    .d(\state[188] ),
    .dl(\state[187] ),
    .dr(\state[189] ),
    .in_data(net4),
    .l(\state[203] ),
    .load_in(_12_),
    .load_out(net114),
    .out_data(\cell_outs[204] ),
    .prev_out_data(\cell_outs[220] ),
    .r(\state[205] ),
    .reset(net70),
    .run(net61),
    .shift(net85),
    .state(\state[204] ),
    .u(\state[220] ),
    .ul(\state[219] ),
    .ur(\state[221] ));
 life_cell arr_cell_x12_y13 (.clk(clknet_5_30__leaf_clk),
    .d(\state[204] ),
    .dl(\state[203] ),
    .dr(\state[205] ),
    .in_data(net4),
    .l(\state[219] ),
    .load_in(_13_),
    .load_out(net114),
    .out_data(\cell_outs[220] ),
    .prev_out_data(\cell_outs[236] ),
    .r(\state[221] ),
    .reset(net70),
    .run(net60),
    .shift(net85),
    .state(\state[220] ),
    .u(\state[236] ),
    .ul(\state[235] ),
    .ur(\state[237] ));
 life_cell arr_cell_x12_y14 (.clk(clknet_5_31__leaf_clk),
    .d(\state[220] ),
    .dl(\state[219] ),
    .dr(\state[221] ),
    .in_data(net4),
    .l(\state[235] ),
    .load_in(_14_),
    .load_out(net114),
    .out_data(\cell_outs[236] ),
    .prev_out_data(\cell_outs[252] ),
    .r(\state[237] ),
    .reset(net70),
    .run(net59),
    .shift(net85),
    .state(\state[236] ),
    .u(\state[252] ),
    .ul(\state[251] ),
    .ur(\state[253] ));
 life_cell arr_cell_x12_y15 (.clk(clknet_5_31__leaf_clk),
    .d(\state[236] ),
    .dl(\state[235] ),
    .dr(\state[237] ),
    .in_data(net4),
    .l(\state[251] ),
    .load_in(_15_),
    .load_out(net114),
    .out_data(\cell_outs[252] ),
    .prev_out_data(net193),
    .r(\state[253] ),
    .reset(net70),
    .run(net58),
    .shift(net85),
    .state(\state[252] ),
    .u(net194),
    .ul(net195),
    .ur(net196));
 life_cell arr_cell_x12_y2 (.clk(clknet_5_11__leaf_clk),
    .d(\state[28] ),
    .dl(\state[27] ),
    .dr(\state[29] ),
    .in_data(net4),
    .l(\state[43] ),
    .load_in(_00_),
    .load_out(net114),
    .out_data(\cell_outs[44] ),
    .prev_out_data(\cell_outs[60] ),
    .r(\state[45] ),
    .reset(net70),
    .run(net54),
    .shift(net85),
    .state(\state[44] ),
    .u(\state[60] ),
    .ul(\state[59] ),
    .ur(\state[61] ));
 life_cell arr_cell_x12_y3 (.clk(clknet_5_11__leaf_clk),
    .d(\state[44] ),
    .dl(\state[43] ),
    .dr(\state[45] ),
    .in_data(net4),
    .l(\state[59] ),
    .load_in(_02_),
    .load_out(net114),
    .out_data(\cell_outs[60] ),
    .prev_out_data(\cell_outs[76] ),
    .r(\state[61] ),
    .reset(net70),
    .run(net55),
    .shift(net85),
    .state(\state[60] ),
    .u(\state[76] ),
    .ul(\state[75] ),
    .ur(\state[77] ));
 life_cell arr_cell_x12_y4 (.clk(clknet_5_14__leaf_clk),
    .d(\state[60] ),
    .dl(\state[59] ),
    .dr(\state[61] ),
    .in_data(net4),
    .l(\state[75] ),
    .load_in(_03_),
    .load_out(net114),
    .out_data(\cell_outs[76] ),
    .prev_out_data(\cell_outs[92] ),
    .r(\state[77] ),
    .reset(net70),
    .run(net56),
    .shift(net85),
    .state(\state[76] ),
    .u(\state[92] ),
    .ul(\state[91] ),
    .ur(\state[93] ));
 life_cell arr_cell_x12_y5 (.clk(clknet_5_14__leaf_clk),
    .d(\state[76] ),
    .dl(\state[75] ),
    .dr(\state[77] ),
    .in_data(net4),
    .l(\state[91] ),
    .load_in(_04_),
    .load_out(net114),
    .out_data(\cell_outs[92] ),
    .prev_out_data(\cell_outs[108] ),
    .r(\state[93] ),
    .reset(net70),
    .run(net57),
    .shift(net85),
    .state(\state[92] ),
    .u(\state[108] ),
    .ul(\state[107] ),
    .ur(\state[109] ));
 life_cell arr_cell_x12_y6 (.clk(clknet_5_15__leaf_clk),
    .d(\state[92] ),
    .dl(\state[91] ),
    .dr(\state[93] ),
    .in_data(net4),
    .l(\state[107] ),
    .load_in(_05_),
    .load_out(net114),
    .out_data(\cell_outs[108] ),
    .prev_out_data(\cell_outs[124] ),
    .r(\state[109] ),
    .reset(net70),
    .run(net66),
    .shift(net85),
    .state(\state[108] ),
    .u(\state[124] ),
    .ul(\state[123] ),
    .ur(\state[125] ));
 life_cell arr_cell_x12_y7 (.clk(clknet_5_15__leaf_clk),
    .d(\state[108] ),
    .dl(\state[107] ),
    .dr(\state[109] ),
    .in_data(net4),
    .l(\state[123] ),
    .load_in(_06_),
    .load_out(net114),
    .out_data(\cell_outs[124] ),
    .prev_out_data(\cell_outs[140] ),
    .r(\state[125] ),
    .reset(net70),
    .run(net25),
    .shift(net85),
    .state(\state[124] ),
    .u(\state[140] ),
    .ul(\state[139] ),
    .ur(\state[141] ));
 life_cell arr_cell_x12_y8 (.clk(clknet_5_26__leaf_clk),
    .d(\state[124] ),
    .dl(\state[123] ),
    .dr(\state[125] ),
    .in_data(net4),
    .l(\state[139] ),
    .load_in(_07_),
    .load_out(net114),
    .out_data(\cell_outs[140] ),
    .prev_out_data(\cell_outs[156] ),
    .r(\state[141] ),
    .reset(net70),
    .run(net65),
    .shift(net85),
    .state(\state[140] ),
    .u(\state[156] ),
    .ul(\state[155] ),
    .ur(\state[157] ));
 life_cell arr_cell_x12_y9 (.clk(clknet_5_26__leaf_clk),
    .d(\state[140] ),
    .dl(\state[139] ),
    .dr(\state[141] ),
    .in_data(net4),
    .l(\state[155] ),
    .load_in(_08_),
    .load_out(net114),
    .out_data(\cell_outs[156] ),
    .prev_out_data(\cell_outs[172] ),
    .r(\state[157] ),
    .reset(net70),
    .run(net64),
    .shift(net85),
    .state(\state[156] ),
    .u(\state[172] ),
    .ul(\state[171] ),
    .ur(\state[173] ));
 life_cell arr_cell_x13_y0 (.clk(clknet_5_10__leaf_clk),
    .d(net197),
    .dl(net198),
    .dr(net199),
    .in_data(net5),
    .l(\state[12] ),
    .load_in(net43),
    .load_out(net113),
    .out_data(\cell_outs[13] ),
    .prev_out_data(\cell_outs[29] ),
    .r(\state[14] ),
    .reset(net69),
    .run(net52),
    .shift(net84),
    .state(\state[13] ),
    .u(\state[29] ),
    .ul(\state[28] ),
    .ur(\state[30] ));
 life_cell arr_cell_x13_y1 (.clk(clknet_5_10__leaf_clk),
    .d(\state[13] ),
    .dl(\state[12] ),
    .dr(\state[14] ),
    .in_data(net5),
    .l(\state[28] ),
    .load_in(_11_),
    .load_out(net113),
    .out_data(\cell_outs[29] ),
    .prev_out_data(\cell_outs[45] ),
    .r(\state[30] ),
    .reset(net69),
    .run(net53),
    .shift(net84),
    .state(\state[29] ),
    .u(\state[45] ),
    .ul(\state[44] ),
    .ur(\state[46] ));
 life_cell arr_cell_x13_y10 (.clk(clknet_5_27__leaf_clk),
    .d(\state[157] ),
    .dl(\state[156] ),
    .dr(\state[158] ),
    .in_data(net5),
    .l(\state[172] ),
    .load_in(_09_),
    .load_out(net113),
    .out_data(\cell_outs[173] ),
    .prev_out_data(\cell_outs[189] ),
    .r(\state[174] ),
    .reset(net69),
    .run(net63),
    .shift(net84),
    .state(\state[173] ),
    .u(\state[189] ),
    .ul(\state[188] ),
    .ur(\state[190] ));
 life_cell arr_cell_x13_y11 (.clk(clknet_5_27__leaf_clk),
    .d(\state[173] ),
    .dl(\state[172] ),
    .dr(\state[174] ),
    .in_data(net5),
    .l(\state[188] ),
    .load_in(_10_),
    .load_out(net113),
    .out_data(\cell_outs[189] ),
    .prev_out_data(\cell_outs[205] ),
    .r(\state[190] ),
    .reset(net69),
    .run(net62),
    .shift(net84),
    .state(\state[189] ),
    .u(\state[205] ),
    .ul(\state[204] ),
    .ur(\state[206] ));
 life_cell arr_cell_x13_y12 (.clk(clknet_5_30__leaf_clk),
    .d(\state[189] ),
    .dl(\state[188] ),
    .dr(\state[190] ),
    .in_data(net5),
    .l(\state[204] ),
    .load_in(_12_),
    .load_out(net113),
    .out_data(\cell_outs[205] ),
    .prev_out_data(\cell_outs[221] ),
    .r(\state[206] ),
    .reset(net69),
    .run(net61),
    .shift(net84),
    .state(\state[205] ),
    .u(\state[221] ),
    .ul(\state[220] ),
    .ur(\state[222] ));
 life_cell arr_cell_x13_y13 (.clk(clknet_5_30__leaf_clk),
    .d(\state[205] ),
    .dl(\state[204] ),
    .dr(\state[206] ),
    .in_data(net5),
    .l(\state[220] ),
    .load_in(_13_),
    .load_out(net113),
    .out_data(\cell_outs[221] ),
    .prev_out_data(\cell_outs[237] ),
    .r(\state[222] ),
    .reset(net69),
    .run(net60),
    .shift(net84),
    .state(\state[221] ),
    .u(\state[237] ),
    .ul(\state[236] ),
    .ur(\state[238] ));
 life_cell arr_cell_x13_y14 (.clk(clknet_5_31__leaf_clk),
    .d(\state[221] ),
    .dl(\state[220] ),
    .dr(\state[222] ),
    .in_data(net5),
    .l(\state[236] ),
    .load_in(_14_),
    .load_out(net113),
    .out_data(\cell_outs[237] ),
    .prev_out_data(\cell_outs[253] ),
    .r(\state[238] ),
    .reset(net69),
    .run(net59),
    .shift(net84),
    .state(\state[237] ),
    .u(\state[253] ),
    .ul(\state[252] ),
    .ur(\state[254] ));
 life_cell arr_cell_x13_y15 (.clk(clknet_5_31__leaf_clk),
    .d(\state[237] ),
    .dl(\state[236] ),
    .dr(\state[238] ),
    .in_data(net5),
    .l(\state[252] ),
    .load_in(_15_),
    .load_out(net113),
    .out_data(\cell_outs[253] ),
    .prev_out_data(net200),
    .r(\state[254] ),
    .reset(net69),
    .run(net58),
    .shift(net84),
    .state(\state[253] ),
    .u(net201),
    .ul(net202),
    .ur(net203));
 life_cell arr_cell_x13_y2 (.clk(clknet_5_11__leaf_clk),
    .d(\state[29] ),
    .dl(\state[28] ),
    .dr(\state[30] ),
    .in_data(net5),
    .l(\state[44] ),
    .load_in(_00_),
    .load_out(net113),
    .out_data(\cell_outs[45] ),
    .prev_out_data(\cell_outs[61] ),
    .r(\state[46] ),
    .reset(net69),
    .run(net54),
    .shift(net84),
    .state(\state[45] ),
    .u(\state[61] ),
    .ul(\state[60] ),
    .ur(\state[62] ));
 life_cell arr_cell_x13_y3 (.clk(clknet_5_11__leaf_clk),
    .d(\state[45] ),
    .dl(\state[44] ),
    .dr(\state[46] ),
    .in_data(net5),
    .l(\state[60] ),
    .load_in(_02_),
    .load_out(net113),
    .out_data(\cell_outs[61] ),
    .prev_out_data(\cell_outs[77] ),
    .r(\state[62] ),
    .reset(net69),
    .run(net55),
    .shift(net84),
    .state(\state[61] ),
    .u(\state[77] ),
    .ul(\state[76] ),
    .ur(\state[78] ));
 life_cell arr_cell_x13_y4 (.clk(clknet_5_14__leaf_clk),
    .d(\state[61] ),
    .dl(\state[60] ),
    .dr(\state[62] ),
    .in_data(net5),
    .l(\state[76] ),
    .load_in(_03_),
    .load_out(net113),
    .out_data(\cell_outs[77] ),
    .prev_out_data(\cell_outs[93] ),
    .r(\state[78] ),
    .reset(net69),
    .run(net56),
    .shift(net84),
    .state(\state[77] ),
    .u(\state[93] ),
    .ul(\state[92] ),
    .ur(\state[94] ));
 life_cell arr_cell_x13_y5 (.clk(clknet_5_14__leaf_clk),
    .d(\state[77] ),
    .dl(\state[76] ),
    .dr(\state[78] ),
    .in_data(net5),
    .l(\state[92] ),
    .load_in(_04_),
    .load_out(net113),
    .out_data(\cell_outs[93] ),
    .prev_out_data(\cell_outs[109] ),
    .r(\state[94] ),
    .reset(net69),
    .run(net57),
    .shift(net84),
    .state(\state[93] ),
    .u(\state[109] ),
    .ul(\state[108] ),
    .ur(\state[110] ));
 life_cell arr_cell_x13_y6 (.clk(clknet_5_15__leaf_clk),
    .d(\state[93] ),
    .dl(\state[92] ),
    .dr(\state[94] ),
    .in_data(net5),
    .l(\state[108] ),
    .load_in(_05_),
    .load_out(net113),
    .out_data(\cell_outs[109] ),
    .prev_out_data(\cell_outs[125] ),
    .r(\state[110] ),
    .reset(net69),
    .run(net66),
    .shift(net84),
    .state(\state[109] ),
    .u(\state[125] ),
    .ul(\state[124] ),
    .ur(\state[126] ));
 life_cell arr_cell_x13_y7 (.clk(clknet_5_15__leaf_clk),
    .d(\state[109] ),
    .dl(\state[108] ),
    .dr(\state[110] ),
    .in_data(net5),
    .l(\state[124] ),
    .load_in(_06_),
    .load_out(net113),
    .out_data(\cell_outs[125] ),
    .prev_out_data(\cell_outs[141] ),
    .r(\state[126] ),
    .reset(net69),
    .run(net25),
    .shift(net84),
    .state(\state[125] ),
    .u(\state[141] ),
    .ul(\state[140] ),
    .ur(\state[142] ));
 life_cell arr_cell_x13_y8 (.clk(clknet_5_26__leaf_clk),
    .d(\state[125] ),
    .dl(\state[124] ),
    .dr(\state[126] ),
    .in_data(net5),
    .l(\state[140] ),
    .load_in(_07_),
    .load_out(net113),
    .out_data(\cell_outs[141] ),
    .prev_out_data(\cell_outs[157] ),
    .r(\state[142] ),
    .reset(net69),
    .run(net65),
    .shift(net84),
    .state(\state[141] ),
    .u(\state[157] ),
    .ul(\state[156] ),
    .ur(\state[158] ));
 life_cell arr_cell_x13_y9 (.clk(clknet_5_26__leaf_clk),
    .d(\state[141] ),
    .dl(\state[140] ),
    .dr(\state[142] ),
    .in_data(net5),
    .l(\state[156] ),
    .load_in(_08_),
    .load_out(net113),
    .out_data(\cell_outs[157] ),
    .prev_out_data(\cell_outs[173] ),
    .r(\state[158] ),
    .reset(net69),
    .run(net64),
    .shift(net84),
    .state(\state[157] ),
    .u(\state[173] ),
    .ul(\state[172] ),
    .ur(\state[174] ));
 life_cell arr_cell_x14_y0 (.clk(clknet_5_10__leaf_clk),
    .d(net204),
    .dl(net205),
    .dr(net206),
    .in_data(net6),
    .l(\state[13] ),
    .load_in(net43),
    .load_out(net112),
    .out_data(\cell_outs[14] ),
    .prev_out_data(\cell_outs[30] ),
    .r(\state[15] ),
    .reset(net68),
    .run(net52),
    .shift(net83),
    .state(\state[14] ),
    .u(\state[30] ),
    .ul(\state[29] ),
    .ur(\state[31] ));
 life_cell arr_cell_x14_y1 (.clk(clknet_5_10__leaf_clk),
    .d(\state[14] ),
    .dl(\state[13] ),
    .dr(\state[15] ),
    .in_data(net6),
    .l(\state[29] ),
    .load_in(_11_),
    .load_out(net112),
    .out_data(\cell_outs[30] ),
    .prev_out_data(\cell_outs[46] ),
    .r(\state[31] ),
    .reset(net68),
    .run(net53),
    .shift(net83),
    .state(\state[30] ),
    .u(\state[46] ),
    .ul(\state[45] ),
    .ur(\state[47] ));
 life_cell arr_cell_x14_y10 (.clk(clknet_5_27__leaf_clk),
    .d(\state[158] ),
    .dl(\state[157] ),
    .dr(\state[159] ),
    .in_data(net6),
    .l(\state[173] ),
    .load_in(_09_),
    .load_out(net112),
    .out_data(\cell_outs[174] ),
    .prev_out_data(\cell_outs[190] ),
    .r(\state[175] ),
    .reset(net68),
    .run(net63),
    .shift(net83),
    .state(\state[174] ),
    .u(\state[190] ),
    .ul(\state[189] ),
    .ur(\state[191] ));
 life_cell arr_cell_x14_y11 (.clk(clknet_5_27__leaf_clk),
    .d(\state[174] ),
    .dl(\state[173] ),
    .dr(\state[175] ),
    .in_data(net6),
    .l(\state[189] ),
    .load_in(_10_),
    .load_out(net112),
    .out_data(\cell_outs[190] ),
    .prev_out_data(\cell_outs[206] ),
    .r(\state[191] ),
    .reset(net68),
    .run(net62),
    .shift(net83),
    .state(\state[190] ),
    .u(\state[206] ),
    .ul(\state[205] ),
    .ur(\state[207] ));
 life_cell arr_cell_x14_y12 (.clk(clknet_5_30__leaf_clk),
    .d(\state[190] ),
    .dl(\state[189] ),
    .dr(\state[191] ),
    .in_data(net6),
    .l(\state[205] ),
    .load_in(_12_),
    .load_out(net112),
    .out_data(\cell_outs[206] ),
    .prev_out_data(\cell_outs[222] ),
    .r(\state[207] ),
    .reset(net68),
    .run(net61),
    .shift(net83),
    .state(\state[206] ),
    .u(\state[222] ),
    .ul(\state[221] ),
    .ur(\state[223] ));
 life_cell arr_cell_x14_y13 (.clk(clknet_5_30__leaf_clk),
    .d(\state[206] ),
    .dl(\state[205] ),
    .dr(\state[207] ),
    .in_data(net6),
    .l(\state[221] ),
    .load_in(_13_),
    .load_out(net112),
    .out_data(\cell_outs[222] ),
    .prev_out_data(\cell_outs[238] ),
    .r(\state[223] ),
    .reset(net68),
    .run(net60),
    .shift(net83),
    .state(\state[222] ),
    .u(\state[238] ),
    .ul(\state[237] ),
    .ur(\state[239] ));
 life_cell arr_cell_x14_y14 (.clk(clknet_5_31__leaf_clk),
    .d(\state[222] ),
    .dl(\state[221] ),
    .dr(\state[223] ),
    .in_data(net6),
    .l(\state[237] ),
    .load_in(_14_),
    .load_out(net112),
    .out_data(\cell_outs[238] ),
    .prev_out_data(\cell_outs[254] ),
    .r(\state[239] ),
    .reset(net68),
    .run(net59),
    .shift(net83),
    .state(\state[238] ),
    .u(\state[254] ),
    .ul(\state[253] ),
    .ur(\state[255] ));
 life_cell arr_cell_x14_y15 (.clk(clknet_5_31__leaf_clk),
    .d(\state[238] ),
    .dl(\state[237] ),
    .dr(\state[239] ),
    .in_data(net6),
    .l(\state[253] ),
    .load_in(_15_),
    .load_out(net112),
    .out_data(\cell_outs[254] ),
    .prev_out_data(net207),
    .r(\state[255] ),
    .reset(net68),
    .run(net58),
    .shift(net83),
    .state(\state[254] ),
    .u(net208),
    .ul(net209),
    .ur(net210));
 life_cell arr_cell_x14_y2 (.clk(clknet_5_11__leaf_clk),
    .d(\state[30] ),
    .dl(\state[29] ),
    .dr(\state[31] ),
    .in_data(net6),
    .l(\state[45] ),
    .load_in(_00_),
    .load_out(net112),
    .out_data(\cell_outs[46] ),
    .prev_out_data(\cell_outs[62] ),
    .r(\state[47] ),
    .reset(net68),
    .run(net54),
    .shift(net83),
    .state(\state[46] ),
    .u(\state[62] ),
    .ul(\state[61] ),
    .ur(\state[63] ));
 life_cell arr_cell_x14_y3 (.clk(clknet_5_11__leaf_clk),
    .d(\state[46] ),
    .dl(\state[45] ),
    .dr(\state[47] ),
    .in_data(net6),
    .l(\state[61] ),
    .load_in(_02_),
    .load_out(net112),
    .out_data(\cell_outs[62] ),
    .prev_out_data(\cell_outs[78] ),
    .r(\state[63] ),
    .reset(net68),
    .run(net55),
    .shift(net83),
    .state(\state[62] ),
    .u(\state[78] ),
    .ul(\state[77] ),
    .ur(\state[79] ));
 life_cell arr_cell_x14_y4 (.clk(clknet_5_14__leaf_clk),
    .d(\state[62] ),
    .dl(\state[61] ),
    .dr(\state[63] ),
    .in_data(net6),
    .l(\state[77] ),
    .load_in(_03_),
    .load_out(net112),
    .out_data(\cell_outs[78] ),
    .prev_out_data(\cell_outs[94] ),
    .r(\state[79] ),
    .reset(net68),
    .run(net56),
    .shift(net83),
    .state(\state[78] ),
    .u(\state[94] ),
    .ul(\state[93] ),
    .ur(\state[95] ));
 life_cell arr_cell_x14_y5 (.clk(clknet_5_14__leaf_clk),
    .d(\state[78] ),
    .dl(\state[77] ),
    .dr(\state[79] ),
    .in_data(net6),
    .l(\state[93] ),
    .load_in(_04_),
    .load_out(net112),
    .out_data(\cell_outs[94] ),
    .prev_out_data(\cell_outs[110] ),
    .r(\state[95] ),
    .reset(net68),
    .run(net57),
    .shift(net83),
    .state(\state[94] ),
    .u(\state[110] ),
    .ul(\state[109] ),
    .ur(\state[111] ));
 life_cell arr_cell_x14_y6 (.clk(clknet_5_15__leaf_clk),
    .d(\state[94] ),
    .dl(\state[93] ),
    .dr(\state[95] ),
    .in_data(net6),
    .l(\state[109] ),
    .load_in(_05_),
    .load_out(net112),
    .out_data(\cell_outs[110] ),
    .prev_out_data(\cell_outs[126] ),
    .r(\state[111] ),
    .reset(net68),
    .run(net66),
    .shift(net83),
    .state(\state[110] ),
    .u(\state[126] ),
    .ul(\state[125] ),
    .ur(\state[127] ));
 life_cell arr_cell_x14_y7 (.clk(clknet_5_15__leaf_clk),
    .d(\state[110] ),
    .dl(\state[109] ),
    .dr(\state[111] ),
    .in_data(net6),
    .l(\state[125] ),
    .load_in(_06_),
    .load_out(net112),
    .out_data(\cell_outs[126] ),
    .prev_out_data(\cell_outs[142] ),
    .r(\state[127] ),
    .reset(net68),
    .run(net25),
    .shift(net83),
    .state(\state[126] ),
    .u(\state[142] ),
    .ul(\state[141] ),
    .ur(\state[143] ));
 life_cell arr_cell_x14_y8 (.clk(clknet_5_26__leaf_clk),
    .d(\state[126] ),
    .dl(\state[125] ),
    .dr(\state[127] ),
    .in_data(net6),
    .l(\state[141] ),
    .load_in(_07_),
    .load_out(net112),
    .out_data(\cell_outs[142] ),
    .prev_out_data(\cell_outs[158] ),
    .r(\state[143] ),
    .reset(net68),
    .run(net65),
    .shift(net83),
    .state(\state[142] ),
    .u(\state[158] ),
    .ul(\state[157] ),
    .ur(\state[159] ));
 life_cell arr_cell_x14_y9 (.clk(clknet_5_26__leaf_clk),
    .d(\state[142] ),
    .dl(\state[141] ),
    .dr(\state[143] ),
    .in_data(net6),
    .l(\state[157] ),
    .load_in(_08_),
    .load_out(net112),
    .out_data(\cell_outs[158] ),
    .prev_out_data(\cell_outs[174] ),
    .r(\state[159] ),
    .reset(net68),
    .run(net64),
    .shift(net83),
    .state(\state[158] ),
    .u(\state[174] ),
    .ul(\state[173] ),
    .ur(\state[175] ));
 life_cell arr_cell_x15_y0 (.clk(clknet_5_10__leaf_clk),
    .d(net211),
    .dl(net212),
    .dr(net213),
    .in_data(net51),
    .l(\state[14] ),
    .load_in(net43),
    .load_out(net111),
    .out_data(\cell_outs[15] ),
    .prev_out_data(\cell_outs[31] ),
    .r(net214),
    .reset(net67),
    .run(net52),
    .shift(net82),
    .state(\state[15] ),
    .u(\state[31] ),
    .ul(\state[30] ),
    .ur(net215));
 life_cell arr_cell_x15_y1 (.clk(clknet_5_10__leaf_clk),
    .d(\state[15] ),
    .dl(\state[14] ),
    .dr(net216),
    .in_data(net51),
    .l(\state[30] ),
    .load_in(_11_),
    .load_out(net111),
    .out_data(\cell_outs[31] ),
    .prev_out_data(\cell_outs[47] ),
    .r(net217),
    .reset(net67),
    .run(net53),
    .shift(net82),
    .state(\state[31] ),
    .u(\state[47] ),
    .ul(\state[46] ),
    .ur(net218));
 life_cell arr_cell_x15_y10 (.clk(clknet_5_27__leaf_clk),
    .d(\state[159] ),
    .dl(\state[158] ),
    .dr(net219),
    .in_data(net51),
    .l(\state[174] ),
    .load_in(_09_),
    .load_out(net111),
    .out_data(\cell_outs[175] ),
    .prev_out_data(\cell_outs[191] ),
    .r(net220),
    .reset(net67),
    .run(net63),
    .shift(net82),
    .state(\state[175] ),
    .u(\state[191] ),
    .ul(\state[190] ),
    .ur(net221));
 life_cell arr_cell_x15_y11 (.clk(clknet_5_27__leaf_clk),
    .d(\state[175] ),
    .dl(\state[174] ),
    .dr(net222),
    .in_data(net51),
    .l(\state[190] ),
    .load_in(_10_),
    .load_out(net111),
    .out_data(\cell_outs[191] ),
    .prev_out_data(\cell_outs[207] ),
    .r(net223),
    .reset(net67),
    .run(net62),
    .shift(net82),
    .state(\state[191] ),
    .u(\state[207] ),
    .ul(\state[206] ),
    .ur(net224));
 life_cell arr_cell_x15_y12 (.clk(clknet_5_30__leaf_clk),
    .d(\state[191] ),
    .dl(\state[190] ),
    .dr(net225),
    .in_data(net51),
    .l(\state[206] ),
    .load_in(_12_),
    .load_out(net111),
    .out_data(\cell_outs[207] ),
    .prev_out_data(\cell_outs[223] ),
    .r(net226),
    .reset(net67),
    .run(net61),
    .shift(net82),
    .state(\state[207] ),
    .u(\state[223] ),
    .ul(\state[222] ),
    .ur(net227));
 life_cell arr_cell_x15_y13 (.clk(clknet_5_30__leaf_clk),
    .d(\state[207] ),
    .dl(\state[206] ),
    .dr(net228),
    .in_data(net51),
    .l(\state[222] ),
    .load_in(_13_),
    .load_out(net111),
    .out_data(\cell_outs[223] ),
    .prev_out_data(\cell_outs[239] ),
    .r(net229),
    .reset(net67),
    .run(net60),
    .shift(net82),
    .state(\state[223] ),
    .u(\state[239] ),
    .ul(\state[238] ),
    .ur(net230));
 life_cell arr_cell_x15_y14 (.clk(clknet_5_31__leaf_clk),
    .d(\state[223] ),
    .dl(\state[222] ),
    .dr(net231),
    .in_data(net51),
    .l(\state[238] ),
    .load_in(_14_),
    .load_out(net111),
    .out_data(\cell_outs[239] ),
    .prev_out_data(\cell_outs[255] ),
    .r(net232),
    .reset(net67),
    .run(net59),
    .shift(net82),
    .state(\state[239] ),
    .u(\state[255] ),
    .ul(\state[254] ),
    .ur(net233));
 life_cell arr_cell_x15_y15 (.clk(clknet_5_31__leaf_clk),
    .d(\state[239] ),
    .dl(\state[238] ),
    .dr(net234),
    .in_data(net51),
    .l(\state[254] ),
    .load_in(_15_),
    .load_out(net111),
    .out_data(\cell_outs[255] ),
    .prev_out_data(net235),
    .r(net236),
    .reset(net67),
    .run(net58),
    .shift(net82),
    .state(\state[255] ),
    .u(net237),
    .ul(net238),
    .ur(net239));
 life_cell arr_cell_x15_y2 (.clk(clknet_5_11__leaf_clk),
    .d(\state[31] ),
    .dl(\state[30] ),
    .dr(net240),
    .in_data(net51),
    .l(\state[46] ),
    .load_in(_00_),
    .load_out(net111),
    .out_data(\cell_outs[47] ),
    .prev_out_data(\cell_outs[63] ),
    .r(net241),
    .reset(net67),
    .run(net54),
    .shift(net82),
    .state(\state[47] ),
    .u(\state[63] ),
    .ul(\state[62] ),
    .ur(net242));
 life_cell arr_cell_x15_y3 (.clk(clknet_5_11__leaf_clk),
    .d(\state[47] ),
    .dl(\state[46] ),
    .dr(net243),
    .in_data(net51),
    .l(\state[62] ),
    .load_in(_02_),
    .load_out(net111),
    .out_data(\cell_outs[63] ),
    .prev_out_data(\cell_outs[79] ),
    .r(net244),
    .reset(net67),
    .run(net55),
    .shift(net82),
    .state(\state[63] ),
    .u(\state[79] ),
    .ul(\state[78] ),
    .ur(net245));
 life_cell arr_cell_x15_y4 (.clk(clknet_5_14__leaf_clk),
    .d(\state[63] ),
    .dl(\state[62] ),
    .dr(net246),
    .in_data(net51),
    .l(\state[78] ),
    .load_in(_03_),
    .load_out(net111),
    .out_data(\cell_outs[79] ),
    .prev_out_data(\cell_outs[95] ),
    .r(net247),
    .reset(net67),
    .run(net56),
    .shift(net82),
    .state(\state[79] ),
    .u(\state[95] ),
    .ul(\state[94] ),
    .ur(net248));
 life_cell arr_cell_x15_y5 (.clk(clknet_5_14__leaf_clk),
    .d(\state[79] ),
    .dl(\state[78] ),
    .dr(net249),
    .in_data(net51),
    .l(\state[94] ),
    .load_in(_04_),
    .load_out(net111),
    .out_data(\cell_outs[95] ),
    .prev_out_data(\cell_outs[111] ),
    .r(net250),
    .reset(net67),
    .run(net57),
    .shift(net82),
    .state(\state[95] ),
    .u(\state[111] ),
    .ul(\state[110] ),
    .ur(net251));
 life_cell arr_cell_x15_y6 (.clk(clknet_5_15__leaf_clk),
    .d(\state[95] ),
    .dl(\state[94] ),
    .dr(net252),
    .in_data(net51),
    .l(\state[110] ),
    .load_in(_05_),
    .load_out(net111),
    .out_data(\cell_outs[111] ),
    .prev_out_data(\cell_outs[127] ),
    .r(net253),
    .reset(net67),
    .run(net66),
    .shift(net82),
    .state(\state[111] ),
    .u(\state[127] ),
    .ul(\state[126] ),
    .ur(net254));
 life_cell arr_cell_x15_y7 (.clk(clknet_5_15__leaf_clk),
    .d(\state[111] ),
    .dl(\state[110] ),
    .dr(net255),
    .in_data(net51),
    .l(\state[126] ),
    .load_in(_06_),
    .load_out(net111),
    .out_data(\cell_outs[127] ),
    .prev_out_data(\cell_outs[143] ),
    .r(net256),
    .reset(net67),
    .run(net25),
    .shift(net82),
    .state(\state[127] ),
    .u(\state[143] ),
    .ul(\state[142] ),
    .ur(net257));
 life_cell arr_cell_x15_y8 (.clk(clknet_5_26__leaf_clk),
    .d(\state[127] ),
    .dl(\state[126] ),
    .dr(net258),
    .in_data(net51),
    .l(\state[142] ),
    .load_in(_07_),
    .load_out(net111),
    .out_data(\cell_outs[143] ),
    .prev_out_data(\cell_outs[159] ),
    .r(net259),
    .reset(net67),
    .run(net65),
    .shift(net82),
    .state(\state[143] ),
    .u(\state[159] ),
    .ul(\state[158] ),
    .ur(net260));
 life_cell arr_cell_x15_y9 (.clk(clknet_5_26__leaf_clk),
    .d(\state[143] ),
    .dl(\state[142] ),
    .dr(net261),
    .in_data(net51),
    .l(\state[158] ),
    .load_in(_08_),
    .load_out(net111),
    .out_data(\cell_outs[159] ),
    .prev_out_data(\cell_outs[175] ),
    .r(net262),
    .reset(net67),
    .run(net64),
    .shift(net82),
    .state(\state[159] ),
    .u(\state[175] ),
    .ul(\state[174] ),
    .ur(net263));
 life_cell arr_cell_x1_y0 (.clk(clknet_5_0__leaf_clk),
    .d(net264),
    .dl(net265),
    .dr(net266),
    .in_data(net8),
    .l(\state[0] ),
    .load_in(net42),
    .load_out(net22),
    .out_data(\cell_outs[1] ),
    .prev_out_data(\cell_outs[17] ),
    .r(\state[2] ),
    .reset(net81),
    .run(net52),
    .shift(net96),
    .state(\state[1] ),
    .u(\state[17] ),
    .ul(\state[16] ),
    .ur(\state[18] ));
 life_cell arr_cell_x1_y1 (.clk(clknet_5_0__leaf_clk),
    .d(\state[1] ),
    .dl(\state[0] ),
    .dr(\state[2] ),
    .in_data(net8),
    .l(\state[16] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[17] ),
    .prev_out_data(\cell_outs[33] ),
    .r(\state[18] ),
    .reset(net81),
    .run(net53),
    .shift(net96),
    .state(\state[17] ),
    .u(\state[33] ),
    .ul(\state[32] ),
    .ur(\state[34] ));
 life_cell arr_cell_x1_y10 (.clk(clknet_5_17__leaf_clk),
    .d(\state[145] ),
    .dl(\state[144] ),
    .dr(\state[146] ),
    .in_data(net8),
    .l(\state[160] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[161] ),
    .prev_out_data(\cell_outs[177] ),
    .r(\state[162] ),
    .reset(net81),
    .run(net63),
    .shift(net96),
    .state(\state[161] ),
    .u(\state[177] ),
    .ul(\state[176] ),
    .ur(\state[178] ));
 life_cell arr_cell_x1_y11 (.clk(clknet_5_17__leaf_clk),
    .d(\state[161] ),
    .dl(\state[160] ),
    .dr(\state[162] ),
    .in_data(net8),
    .l(\state[176] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[177] ),
    .prev_out_data(\cell_outs[193] ),
    .r(\state[178] ),
    .reset(net81),
    .run(net62),
    .shift(net96),
    .state(\state[177] ),
    .u(\state[193] ),
    .ul(\state[192] ),
    .ur(\state[194] ));
 life_cell arr_cell_x1_y12 (.clk(clknet_5_20__leaf_clk),
    .d(\state[177] ),
    .dl(\state[176] ),
    .dr(\state[178] ),
    .in_data(net8),
    .l(\state[192] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[193] ),
    .prev_out_data(\cell_outs[209] ),
    .r(\state[194] ),
    .reset(net81),
    .run(net61),
    .shift(net96),
    .state(\state[193] ),
    .u(\state[209] ),
    .ul(\state[208] ),
    .ur(\state[210] ));
 life_cell arr_cell_x1_y13 (.clk(clknet_5_20__leaf_clk),
    .d(\state[193] ),
    .dl(\state[192] ),
    .dr(\state[194] ),
    .in_data(net8),
    .l(\state[208] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[209] ),
    .prev_out_data(\cell_outs[225] ),
    .r(\state[210] ),
    .reset(net81),
    .run(net60),
    .shift(net96),
    .state(\state[209] ),
    .u(\state[225] ),
    .ul(\state[224] ),
    .ur(\state[226] ));
 life_cell arr_cell_x1_y14 (.clk(clknet_5_21__leaf_clk),
    .d(\state[209] ),
    .dl(\state[208] ),
    .dr(\state[210] ),
    .in_data(net8),
    .l(\state[224] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[225] ),
    .prev_out_data(\cell_outs[241] ),
    .r(\state[226] ),
    .reset(net81),
    .run(net59),
    .shift(net96),
    .state(\state[225] ),
    .u(\state[241] ),
    .ul(\state[240] ),
    .ur(\state[242] ));
 life_cell arr_cell_x1_y15 (.clk(clknet_5_21__leaf_clk),
    .d(\state[225] ),
    .dl(\state[224] ),
    .dr(\state[226] ),
    .in_data(net8),
    .l(\state[240] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[241] ),
    .prev_out_data(net267),
    .r(\state[242] ),
    .reset(net81),
    .run(net58),
    .shift(net96),
    .state(\state[241] ),
    .u(net268),
    .ul(net269),
    .ur(net270));
 life_cell arr_cell_x1_y2 (.clk(clknet_5_1__leaf_clk),
    .d(\state[17] ),
    .dl(\state[16] ),
    .dr(\state[18] ),
    .in_data(net8),
    .l(\state[32] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[33] ),
    .prev_out_data(\cell_outs[49] ),
    .r(\state[34] ),
    .reset(net81),
    .run(net54),
    .shift(net96),
    .state(\state[33] ),
    .u(\state[49] ),
    .ul(\state[48] ),
    .ur(\state[50] ));
 life_cell arr_cell_x1_y3 (.clk(clknet_5_1__leaf_clk),
    .d(\state[33] ),
    .dl(\state[32] ),
    .dr(\state[34] ),
    .in_data(net8),
    .l(\state[48] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[49] ),
    .prev_out_data(\cell_outs[65] ),
    .r(\state[50] ),
    .reset(net81),
    .run(net55),
    .shift(net96),
    .state(\state[49] ),
    .u(\state[65] ),
    .ul(\state[64] ),
    .ur(\state[66] ));
 life_cell arr_cell_x1_y4 (.clk(clknet_5_4__leaf_clk),
    .d(\state[49] ),
    .dl(\state[48] ),
    .dr(\state[50] ),
    .in_data(net8),
    .l(\state[64] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[65] ),
    .prev_out_data(\cell_outs[81] ),
    .r(\state[66] ),
    .reset(net81),
    .run(net56),
    .shift(net96),
    .state(\state[65] ),
    .u(\state[81] ),
    .ul(\state[80] ),
    .ur(\state[82] ));
 life_cell arr_cell_x1_y5 (.clk(clknet_5_4__leaf_clk),
    .d(\state[65] ),
    .dl(\state[64] ),
    .dr(\state[66] ),
    .in_data(net8),
    .l(\state[80] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[81] ),
    .prev_out_data(\cell_outs[97] ),
    .r(\state[82] ),
    .reset(net81),
    .run(net57),
    .shift(net96),
    .state(\state[81] ),
    .u(\state[97] ),
    .ul(\state[96] ),
    .ur(\state[98] ));
 life_cell arr_cell_x1_y6 (.clk(clknet_5_5__leaf_clk),
    .d(\state[81] ),
    .dl(\state[80] ),
    .dr(\state[82] ),
    .in_data(net8),
    .l(\state[96] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[97] ),
    .prev_out_data(\cell_outs[113] ),
    .r(\state[98] ),
    .reset(net81),
    .run(net66),
    .shift(net96),
    .state(\state[97] ),
    .u(\state[113] ),
    .ul(\state[112] ),
    .ur(\state[114] ));
 life_cell arr_cell_x1_y7 (.clk(clknet_5_5__leaf_clk),
    .d(\state[97] ),
    .dl(\state[96] ),
    .dr(\state[98] ),
    .in_data(net8),
    .l(\state[112] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[113] ),
    .prev_out_data(\cell_outs[129] ),
    .r(\state[114] ),
    .reset(net81),
    .run(net25),
    .shift(net96),
    .state(\state[113] ),
    .u(\state[129] ),
    .ul(\state[128] ),
    .ur(\state[130] ));
 life_cell arr_cell_x1_y8 (.clk(clknet_5_16__leaf_clk),
    .d(\state[113] ),
    .dl(\state[112] ),
    .dr(\state[114] ),
    .in_data(net8),
    .l(\state[128] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[129] ),
    .prev_out_data(\cell_outs[145] ),
    .r(\state[130] ),
    .reset(net81),
    .run(net65),
    .shift(net96),
    .state(\state[129] ),
    .u(\state[145] ),
    .ul(\state[144] ),
    .ur(\state[146] ));
 life_cell arr_cell_x1_y9 (.clk(clknet_5_16__leaf_clk),
    .d(\state[129] ),
    .dl(\state[128] ),
    .dr(\state[130] ),
    .in_data(net8),
    .l(\state[144] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[145] ),
    .prev_out_data(\cell_outs[161] ),
    .r(\state[146] ),
    .reset(net81),
    .run(net64),
    .shift(net96),
    .state(\state[145] ),
    .u(\state[161] ),
    .ul(\state[160] ),
    .ur(\state[162] ));
 life_cell arr_cell_x2_y0 (.clk(clknet_5_0__leaf_clk),
    .d(net271),
    .dl(net272),
    .dr(net273),
    .in_data(net50),
    .l(\state[1] ),
    .load_in(net42),
    .load_out(net22),
    .out_data(\cell_outs[2] ),
    .prev_out_data(\cell_outs[18] ),
    .r(\state[3] ),
    .reset(net80),
    .run(net52),
    .shift(net95),
    .state(\state[2] ),
    .u(\state[18] ),
    .ul(\state[17] ),
    .ur(\state[19] ));
 life_cell arr_cell_x2_y1 (.clk(clknet_5_0__leaf_clk),
    .d(\state[2] ),
    .dl(\state[1] ),
    .dr(\state[3] ),
    .in_data(net50),
    .l(\state[17] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[18] ),
    .prev_out_data(\cell_outs[34] ),
    .r(\state[19] ),
    .reset(net80),
    .run(net53),
    .shift(net95),
    .state(\state[18] ),
    .u(\state[34] ),
    .ul(\state[33] ),
    .ur(\state[35] ));
 life_cell arr_cell_x2_y10 (.clk(clknet_5_17__leaf_clk),
    .d(\state[146] ),
    .dl(\state[145] ),
    .dr(\state[147] ),
    .in_data(net50),
    .l(\state[161] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[162] ),
    .prev_out_data(\cell_outs[178] ),
    .r(\state[163] ),
    .reset(net80),
    .run(net63),
    .shift(net95),
    .state(\state[162] ),
    .u(\state[178] ),
    .ul(\state[177] ),
    .ur(\state[179] ));
 life_cell arr_cell_x2_y11 (.clk(clknet_5_17__leaf_clk),
    .d(\state[162] ),
    .dl(\state[161] ),
    .dr(\state[163] ),
    .in_data(net50),
    .l(\state[177] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[178] ),
    .prev_out_data(\cell_outs[194] ),
    .r(\state[179] ),
    .reset(net80),
    .run(net62),
    .shift(net95),
    .state(\state[178] ),
    .u(\state[194] ),
    .ul(\state[193] ),
    .ur(\state[195] ));
 life_cell arr_cell_x2_y12 (.clk(clknet_5_20__leaf_clk),
    .d(\state[178] ),
    .dl(\state[177] ),
    .dr(\state[179] ),
    .in_data(net50),
    .l(\state[193] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[194] ),
    .prev_out_data(\cell_outs[210] ),
    .r(\state[195] ),
    .reset(net80),
    .run(net61),
    .shift(net95),
    .state(\state[194] ),
    .u(\state[210] ),
    .ul(\state[209] ),
    .ur(\state[211] ));
 life_cell arr_cell_x2_y13 (.clk(clknet_5_20__leaf_clk),
    .d(\state[194] ),
    .dl(\state[193] ),
    .dr(\state[195] ),
    .in_data(net50),
    .l(\state[209] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[210] ),
    .prev_out_data(\cell_outs[226] ),
    .r(\state[211] ),
    .reset(net80),
    .run(net60),
    .shift(net95),
    .state(\state[210] ),
    .u(\state[226] ),
    .ul(\state[225] ),
    .ur(\state[227] ));
 life_cell arr_cell_x2_y14 (.clk(clknet_5_21__leaf_clk),
    .d(\state[210] ),
    .dl(\state[209] ),
    .dr(\state[211] ),
    .in_data(net50),
    .l(\state[225] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[226] ),
    .prev_out_data(\cell_outs[242] ),
    .r(\state[227] ),
    .reset(net80),
    .run(net59),
    .shift(net95),
    .state(\state[226] ),
    .u(\state[242] ),
    .ul(\state[241] ),
    .ur(\state[243] ));
 life_cell arr_cell_x2_y15 (.clk(clknet_5_21__leaf_clk),
    .d(\state[226] ),
    .dl(\state[225] ),
    .dr(\state[227] ),
    .in_data(net50),
    .l(\state[241] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[242] ),
    .prev_out_data(net274),
    .r(\state[243] ),
    .reset(net80),
    .run(net58),
    .shift(net95),
    .state(\state[242] ),
    .u(net275),
    .ul(net276),
    .ur(net277));
 life_cell arr_cell_x2_y2 (.clk(clknet_5_1__leaf_clk),
    .d(\state[18] ),
    .dl(\state[17] ),
    .dr(\state[19] ),
    .in_data(net50),
    .l(\state[33] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[34] ),
    .prev_out_data(\cell_outs[50] ),
    .r(\state[35] ),
    .reset(net80),
    .run(net54),
    .shift(net95),
    .state(\state[34] ),
    .u(\state[50] ),
    .ul(\state[49] ),
    .ur(\state[51] ));
 life_cell arr_cell_x2_y3 (.clk(clknet_5_1__leaf_clk),
    .d(\state[34] ),
    .dl(\state[33] ),
    .dr(\state[35] ),
    .in_data(net50),
    .l(\state[49] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[50] ),
    .prev_out_data(\cell_outs[66] ),
    .r(\state[51] ),
    .reset(net80),
    .run(net55),
    .shift(net95),
    .state(\state[50] ),
    .u(\state[66] ),
    .ul(\state[65] ),
    .ur(\state[67] ));
 life_cell arr_cell_x2_y4 (.clk(clknet_5_4__leaf_clk),
    .d(\state[50] ),
    .dl(\state[49] ),
    .dr(\state[51] ),
    .in_data(net50),
    .l(\state[65] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[66] ),
    .prev_out_data(\cell_outs[82] ),
    .r(\state[67] ),
    .reset(net80),
    .run(net56),
    .shift(net95),
    .state(\state[66] ),
    .u(\state[82] ),
    .ul(\state[81] ),
    .ur(\state[83] ));
 life_cell arr_cell_x2_y5 (.clk(clknet_5_4__leaf_clk),
    .d(\state[66] ),
    .dl(\state[65] ),
    .dr(\state[67] ),
    .in_data(net50),
    .l(\state[81] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[82] ),
    .prev_out_data(\cell_outs[98] ),
    .r(\state[83] ),
    .reset(net80),
    .run(net57),
    .shift(net95),
    .state(\state[82] ),
    .u(\state[98] ),
    .ul(\state[97] ),
    .ur(\state[99] ));
 life_cell arr_cell_x2_y6 (.clk(clknet_5_5__leaf_clk),
    .d(\state[82] ),
    .dl(\state[81] ),
    .dr(\state[83] ),
    .in_data(net50),
    .l(\state[97] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[98] ),
    .prev_out_data(\cell_outs[114] ),
    .r(\state[99] ),
    .reset(net80),
    .run(net66),
    .shift(net95),
    .state(\state[98] ),
    .u(\state[114] ),
    .ul(\state[113] ),
    .ur(\state[115] ));
 life_cell arr_cell_x2_y7 (.clk(clknet_5_5__leaf_clk),
    .d(\state[98] ),
    .dl(\state[97] ),
    .dr(\state[99] ),
    .in_data(net50),
    .l(\state[113] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[114] ),
    .prev_out_data(\cell_outs[130] ),
    .r(\state[115] ),
    .reset(net80),
    .run(net25),
    .shift(net95),
    .state(\state[114] ),
    .u(\state[130] ),
    .ul(\state[129] ),
    .ur(\state[131] ));
 life_cell arr_cell_x2_y8 (.clk(clknet_5_16__leaf_clk),
    .d(\state[114] ),
    .dl(\state[113] ),
    .dr(\state[115] ),
    .in_data(net50),
    .l(\state[129] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[130] ),
    .prev_out_data(\cell_outs[146] ),
    .r(\state[131] ),
    .reset(net80),
    .run(net65),
    .shift(net95),
    .state(\state[130] ),
    .u(\state[146] ),
    .ul(\state[145] ),
    .ur(\state[147] ));
 life_cell arr_cell_x2_y9 (.clk(clknet_5_16__leaf_clk),
    .d(\state[130] ),
    .dl(\state[129] ),
    .dr(\state[131] ),
    .in_data(net50),
    .l(\state[145] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[146] ),
    .prev_out_data(\cell_outs[162] ),
    .r(\state[147] ),
    .reset(net80),
    .run(net64),
    .shift(net95),
    .state(\state[146] ),
    .u(\state[162] ),
    .ul(\state[161] ),
    .ur(\state[163] ));
 life_cell arr_cell_x3_y0 (.clk(clknet_5_0__leaf_clk),
    .d(net278),
    .dl(net279),
    .dr(net280),
    .in_data(net10),
    .l(\state[2] ),
    .load_in(net47),
    .load_out(net22),
    .out_data(\cell_outs[3] ),
    .prev_out_data(\cell_outs[19] ),
    .r(\state[4] ),
    .reset(net79),
    .run(net52),
    .shift(net94),
    .state(\state[3] ),
    .u(\state[19] ),
    .ul(\state[18] ),
    .ur(\state[20] ));
 life_cell arr_cell_x3_y1 (.clk(clknet_5_0__leaf_clk),
    .d(\state[3] ),
    .dl(\state[2] ),
    .dr(\state[4] ),
    .in_data(net10),
    .l(\state[18] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[19] ),
    .prev_out_data(\cell_outs[35] ),
    .r(\state[20] ),
    .reset(net79),
    .run(net53),
    .shift(net94),
    .state(\state[19] ),
    .u(\state[35] ),
    .ul(\state[34] ),
    .ur(\state[36] ));
 life_cell arr_cell_x3_y10 (.clk(clknet_5_17__leaf_clk),
    .d(\state[147] ),
    .dl(\state[146] ),
    .dr(\state[148] ),
    .in_data(net10),
    .l(\state[162] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[163] ),
    .prev_out_data(\cell_outs[179] ),
    .r(\state[164] ),
    .reset(net79),
    .run(net63),
    .shift(net94),
    .state(\state[163] ),
    .u(\state[179] ),
    .ul(\state[178] ),
    .ur(\state[180] ));
 life_cell arr_cell_x3_y11 (.clk(clknet_5_17__leaf_clk),
    .d(\state[163] ),
    .dl(\state[162] ),
    .dr(\state[164] ),
    .in_data(net10),
    .l(\state[178] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[179] ),
    .prev_out_data(\cell_outs[195] ),
    .r(\state[180] ),
    .reset(net79),
    .run(net62),
    .shift(net94),
    .state(\state[179] ),
    .u(\state[195] ),
    .ul(\state[194] ),
    .ur(\state[196] ));
 life_cell arr_cell_x3_y12 (.clk(clknet_5_20__leaf_clk),
    .d(\state[179] ),
    .dl(\state[178] ),
    .dr(\state[180] ),
    .in_data(net10),
    .l(\state[194] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[195] ),
    .prev_out_data(\cell_outs[211] ),
    .r(\state[196] ),
    .reset(net79),
    .run(net61),
    .shift(net94),
    .state(\state[195] ),
    .u(\state[211] ),
    .ul(\state[210] ),
    .ur(\state[212] ));
 life_cell arr_cell_x3_y13 (.clk(clknet_5_20__leaf_clk),
    .d(\state[195] ),
    .dl(\state[194] ),
    .dr(\state[196] ),
    .in_data(net10),
    .l(\state[210] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[211] ),
    .prev_out_data(\cell_outs[227] ),
    .r(\state[212] ),
    .reset(net79),
    .run(net60),
    .shift(net94),
    .state(\state[211] ),
    .u(\state[227] ),
    .ul(\state[226] ),
    .ur(\state[228] ));
 life_cell arr_cell_x3_y14 (.clk(clknet_5_21__leaf_clk),
    .d(\state[211] ),
    .dl(\state[210] ),
    .dr(\state[212] ),
    .in_data(net10),
    .l(\state[226] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[227] ),
    .prev_out_data(\cell_outs[243] ),
    .r(\state[228] ),
    .reset(net79),
    .run(net59),
    .shift(net94),
    .state(\state[227] ),
    .u(\state[243] ),
    .ul(\state[242] ),
    .ur(\state[244] ));
 life_cell arr_cell_x3_y15 (.clk(clknet_5_21__leaf_clk),
    .d(\state[227] ),
    .dl(\state[226] ),
    .dr(\state[228] ),
    .in_data(net10),
    .l(\state[242] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[243] ),
    .prev_out_data(net281),
    .r(\state[244] ),
    .reset(net79),
    .run(net58),
    .shift(net94),
    .state(\state[243] ),
    .u(net282),
    .ul(net283),
    .ur(net284));
 life_cell arr_cell_x3_y2 (.clk(clknet_5_1__leaf_clk),
    .d(\state[19] ),
    .dl(\state[18] ),
    .dr(\state[20] ),
    .in_data(net10),
    .l(\state[34] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[35] ),
    .prev_out_data(\cell_outs[51] ),
    .r(\state[36] ),
    .reset(net79),
    .run(net54),
    .shift(net94),
    .state(\state[35] ),
    .u(\state[51] ),
    .ul(\state[50] ),
    .ur(\state[52] ));
 life_cell arr_cell_x3_y3 (.clk(clknet_5_1__leaf_clk),
    .d(\state[35] ),
    .dl(\state[34] ),
    .dr(\state[36] ),
    .in_data(net10),
    .l(\state[50] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[51] ),
    .prev_out_data(\cell_outs[67] ),
    .r(\state[52] ),
    .reset(net79),
    .run(net55),
    .shift(net94),
    .state(\state[51] ),
    .u(\state[67] ),
    .ul(\state[66] ),
    .ur(\state[68] ));
 life_cell arr_cell_x3_y4 (.clk(clknet_5_4__leaf_clk),
    .d(\state[51] ),
    .dl(\state[50] ),
    .dr(\state[52] ),
    .in_data(net10),
    .l(\state[66] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[67] ),
    .prev_out_data(\cell_outs[83] ),
    .r(\state[68] ),
    .reset(net79),
    .run(net56),
    .shift(net94),
    .state(\state[67] ),
    .u(\state[83] ),
    .ul(\state[82] ),
    .ur(\state[84] ));
 life_cell arr_cell_x3_y5 (.clk(clknet_5_4__leaf_clk),
    .d(\state[67] ),
    .dl(\state[66] ),
    .dr(\state[68] ),
    .in_data(net10),
    .l(\state[82] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[83] ),
    .prev_out_data(\cell_outs[99] ),
    .r(\state[84] ),
    .reset(net79),
    .run(net57),
    .shift(net94),
    .state(\state[83] ),
    .u(\state[99] ),
    .ul(\state[98] ),
    .ur(\state[100] ));
 life_cell arr_cell_x3_y6 (.clk(clknet_5_5__leaf_clk),
    .d(\state[83] ),
    .dl(\state[82] ),
    .dr(\state[84] ),
    .in_data(net10),
    .l(\state[98] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[99] ),
    .prev_out_data(\cell_outs[115] ),
    .r(\state[100] ),
    .reset(net79),
    .run(net66),
    .shift(net94),
    .state(\state[99] ),
    .u(\state[115] ),
    .ul(\state[114] ),
    .ur(\state[116] ));
 life_cell arr_cell_x3_y7 (.clk(clknet_5_5__leaf_clk),
    .d(\state[99] ),
    .dl(\state[98] ),
    .dr(\state[100] ),
    .in_data(net10),
    .l(\state[114] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[115] ),
    .prev_out_data(\cell_outs[131] ),
    .r(\state[116] ),
    .reset(net79),
    .run(net25),
    .shift(net94),
    .state(\state[115] ),
    .u(\state[131] ),
    .ul(\state[130] ),
    .ur(\state[132] ));
 life_cell arr_cell_x3_y8 (.clk(clknet_5_16__leaf_clk),
    .d(\state[115] ),
    .dl(\state[114] ),
    .dr(\state[116] ),
    .in_data(net10),
    .l(\state[130] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[131] ),
    .prev_out_data(\cell_outs[147] ),
    .r(\state[132] ),
    .reset(net79),
    .run(net65),
    .shift(net94),
    .state(\state[131] ),
    .u(\state[147] ),
    .ul(\state[146] ),
    .ur(\state[148] ));
 life_cell arr_cell_x3_y9 (.clk(clknet_5_16__leaf_clk),
    .d(\state[131] ),
    .dl(\state[130] ),
    .dr(\state[132] ),
    .in_data(net10),
    .l(\state[146] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[147] ),
    .prev_out_data(\cell_outs[163] ),
    .r(\state[148] ),
    .reset(net79),
    .run(net64),
    .shift(net94),
    .state(\state[147] ),
    .u(\state[163] ),
    .ul(\state[162] ),
    .ur(\state[164] ));
 life_cell arr_cell_x4_y0 (.clk(clknet_5_2__leaf_clk),
    .d(net285),
    .dl(net286),
    .dr(net287),
    .in_data(net11),
    .l(\state[3] ),
    .load_in(net47),
    .load_out(net22),
    .out_data(\cell_outs[4] ),
    .prev_out_data(\cell_outs[20] ),
    .r(\state[5] ),
    .reset(net78),
    .run(net52),
    .shift(net93),
    .state(\state[4] ),
    .u(\state[20] ),
    .ul(\state[19] ),
    .ur(\state[21] ));
 life_cell arr_cell_x4_y1 (.clk(clknet_5_2__leaf_clk),
    .d(\state[4] ),
    .dl(\state[3] ),
    .dr(\state[5] ),
    .in_data(net11),
    .l(\state[19] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[20] ),
    .prev_out_data(\cell_outs[36] ),
    .r(\state[21] ),
    .reset(net78),
    .run(net53),
    .shift(net93),
    .state(\state[20] ),
    .u(\state[36] ),
    .ul(\state[35] ),
    .ur(\state[37] ));
 life_cell arr_cell_x4_y10 (.clk(clknet_5_19__leaf_clk),
    .d(\state[148] ),
    .dl(\state[147] ),
    .dr(\state[149] ),
    .in_data(net11),
    .l(\state[163] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[164] ),
    .prev_out_data(\cell_outs[180] ),
    .r(\state[165] ),
    .reset(net78),
    .run(net63),
    .shift(net93),
    .state(\state[164] ),
    .u(\state[180] ),
    .ul(\state[179] ),
    .ur(\state[181] ));
 life_cell arr_cell_x4_y11 (.clk(clknet_5_19__leaf_clk),
    .d(\state[164] ),
    .dl(\state[163] ),
    .dr(\state[165] ),
    .in_data(net11),
    .l(\state[179] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[180] ),
    .prev_out_data(\cell_outs[196] ),
    .r(\state[181] ),
    .reset(net78),
    .run(net62),
    .shift(net93),
    .state(\state[180] ),
    .u(\state[196] ),
    .ul(\state[195] ),
    .ur(\state[197] ));
 life_cell arr_cell_x4_y12 (.clk(clknet_5_22__leaf_clk),
    .d(\state[180] ),
    .dl(\state[179] ),
    .dr(\state[181] ),
    .in_data(net11),
    .l(\state[195] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[196] ),
    .prev_out_data(\cell_outs[212] ),
    .r(\state[197] ),
    .reset(net78),
    .run(net61),
    .shift(net93),
    .state(\state[196] ),
    .u(\state[212] ),
    .ul(\state[211] ),
    .ur(\state[213] ));
 life_cell arr_cell_x4_y13 (.clk(clknet_5_22__leaf_clk),
    .d(\state[196] ),
    .dl(\state[195] ),
    .dr(\state[197] ),
    .in_data(net11),
    .l(\state[211] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[212] ),
    .prev_out_data(\cell_outs[228] ),
    .r(\state[213] ),
    .reset(net78),
    .run(net60),
    .shift(net93),
    .state(\state[212] ),
    .u(\state[228] ),
    .ul(\state[227] ),
    .ur(\state[229] ));
 life_cell arr_cell_x4_y14 (.clk(clknet_5_23__leaf_clk),
    .d(\state[212] ),
    .dl(\state[211] ),
    .dr(\state[213] ),
    .in_data(net11),
    .l(\state[227] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[228] ),
    .prev_out_data(\cell_outs[244] ),
    .r(\state[229] ),
    .reset(net78),
    .run(net59),
    .shift(net93),
    .state(\state[228] ),
    .u(\state[244] ),
    .ul(\state[243] ),
    .ur(\state[245] ));
 life_cell arr_cell_x4_y15 (.clk(clknet_5_23__leaf_clk),
    .d(\state[228] ),
    .dl(\state[227] ),
    .dr(\state[229] ),
    .in_data(net11),
    .l(\state[243] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[244] ),
    .prev_out_data(net288),
    .r(\state[245] ),
    .reset(net78),
    .run(net58),
    .shift(net93),
    .state(\state[244] ),
    .u(net289),
    .ul(net290),
    .ur(net291));
 life_cell arr_cell_x4_y2 (.clk(clknet_5_3__leaf_clk),
    .d(\state[20] ),
    .dl(\state[19] ),
    .dr(\state[21] ),
    .in_data(net11),
    .l(\state[35] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[36] ),
    .prev_out_data(\cell_outs[52] ),
    .r(\state[37] ),
    .reset(net78),
    .run(net54),
    .shift(net93),
    .state(\state[36] ),
    .u(\state[52] ),
    .ul(\state[51] ),
    .ur(\state[53] ));
 life_cell arr_cell_x4_y3 (.clk(clknet_5_3__leaf_clk),
    .d(\state[36] ),
    .dl(\state[35] ),
    .dr(\state[37] ),
    .in_data(net11),
    .l(\state[51] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[52] ),
    .prev_out_data(\cell_outs[68] ),
    .r(\state[53] ),
    .reset(net78),
    .run(net55),
    .shift(net93),
    .state(\state[52] ),
    .u(\state[68] ),
    .ul(\state[67] ),
    .ur(\state[69] ));
 life_cell arr_cell_x4_y4 (.clk(clknet_5_6__leaf_clk),
    .d(\state[52] ),
    .dl(\state[51] ),
    .dr(\state[53] ),
    .in_data(net11),
    .l(\state[67] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[68] ),
    .prev_out_data(\cell_outs[84] ),
    .r(\state[69] ),
    .reset(net78),
    .run(net56),
    .shift(net93),
    .state(\state[68] ),
    .u(\state[84] ),
    .ul(\state[83] ),
    .ur(\state[85] ));
 life_cell arr_cell_x4_y5 (.clk(clknet_5_6__leaf_clk),
    .d(\state[68] ),
    .dl(\state[67] ),
    .dr(\state[69] ),
    .in_data(net11),
    .l(\state[83] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[84] ),
    .prev_out_data(\cell_outs[100] ),
    .r(\state[85] ),
    .reset(net78),
    .run(net57),
    .shift(net93),
    .state(\state[84] ),
    .u(\state[100] ),
    .ul(\state[99] ),
    .ur(\state[101] ));
 life_cell arr_cell_x4_y6 (.clk(clknet_5_7__leaf_clk),
    .d(\state[84] ),
    .dl(\state[83] ),
    .dr(\state[85] ),
    .in_data(net11),
    .l(\state[99] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[100] ),
    .prev_out_data(\cell_outs[116] ),
    .r(\state[101] ),
    .reset(net78),
    .run(net66),
    .shift(net93),
    .state(\state[100] ),
    .u(\state[116] ),
    .ul(\state[115] ),
    .ur(\state[117] ));
 life_cell arr_cell_x4_y7 (.clk(clknet_5_7__leaf_clk),
    .d(\state[100] ),
    .dl(\state[99] ),
    .dr(\state[101] ),
    .in_data(net11),
    .l(\state[115] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[116] ),
    .prev_out_data(\cell_outs[132] ),
    .r(\state[117] ),
    .reset(net78),
    .run(net25),
    .shift(net93),
    .state(\state[116] ),
    .u(\state[132] ),
    .ul(\state[131] ),
    .ur(\state[133] ));
 life_cell arr_cell_x4_y8 (.clk(clknet_5_18__leaf_clk),
    .d(\state[116] ),
    .dl(\state[115] ),
    .dr(\state[117] ),
    .in_data(net11),
    .l(\state[131] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[132] ),
    .prev_out_data(\cell_outs[148] ),
    .r(\state[133] ),
    .reset(net78),
    .run(net65),
    .shift(net93),
    .state(\state[132] ),
    .u(\state[148] ),
    .ul(\state[147] ),
    .ur(\state[149] ));
 life_cell arr_cell_x4_y9 (.clk(clknet_5_18__leaf_clk),
    .d(\state[132] ),
    .dl(\state[131] ),
    .dr(\state[133] ),
    .in_data(net11),
    .l(\state[147] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[148] ),
    .prev_out_data(\cell_outs[164] ),
    .r(\state[149] ),
    .reset(net78),
    .run(net64),
    .shift(net93),
    .state(\state[148] ),
    .u(\state[164] ),
    .ul(\state[163] ),
    .ur(\state[165] ));
 life_cell arr_cell_x5_y0 (.clk(clknet_5_2__leaf_clk),
    .d(net292),
    .dl(net293),
    .dr(net294),
    .in_data(net12),
    .l(\state[4] ),
    .load_in(net47),
    .load_out(net22),
    .out_data(\cell_outs[5] ),
    .prev_out_data(\cell_outs[21] ),
    .r(\state[6] ),
    .reset(net77),
    .run(net52),
    .shift(net92),
    .state(\state[5] ),
    .u(\state[21] ),
    .ul(\state[20] ),
    .ur(\state[22] ));
 life_cell arr_cell_x5_y1 (.clk(clknet_5_2__leaf_clk),
    .d(\state[5] ),
    .dl(\state[4] ),
    .dr(\state[6] ),
    .in_data(net12),
    .l(\state[20] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[21] ),
    .prev_out_data(\cell_outs[37] ),
    .r(\state[22] ),
    .reset(net77),
    .run(net53),
    .shift(net92),
    .state(\state[21] ),
    .u(\state[37] ),
    .ul(\state[36] ),
    .ur(\state[38] ));
 life_cell arr_cell_x5_y10 (.clk(clknet_5_19__leaf_clk),
    .d(\state[149] ),
    .dl(\state[148] ),
    .dr(\state[150] ),
    .in_data(net12),
    .l(\state[164] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[165] ),
    .prev_out_data(\cell_outs[181] ),
    .r(\state[166] ),
    .reset(net77),
    .run(net63),
    .shift(net92),
    .state(\state[165] ),
    .u(\state[181] ),
    .ul(\state[180] ),
    .ur(\state[182] ));
 life_cell arr_cell_x5_y11 (.clk(clknet_5_19__leaf_clk),
    .d(\state[165] ),
    .dl(\state[164] ),
    .dr(\state[166] ),
    .in_data(net12),
    .l(\state[180] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[181] ),
    .prev_out_data(\cell_outs[197] ),
    .r(\state[182] ),
    .reset(net77),
    .run(net62),
    .shift(net92),
    .state(\state[181] ),
    .u(\state[197] ),
    .ul(\state[196] ),
    .ur(\state[198] ));
 life_cell arr_cell_x5_y12 (.clk(clknet_5_22__leaf_clk),
    .d(\state[181] ),
    .dl(\state[180] ),
    .dr(\state[182] ),
    .in_data(net12),
    .l(\state[196] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[197] ),
    .prev_out_data(\cell_outs[213] ),
    .r(\state[198] ),
    .reset(net77),
    .run(net61),
    .shift(net92),
    .state(\state[197] ),
    .u(\state[213] ),
    .ul(\state[212] ),
    .ur(\state[214] ));
 life_cell arr_cell_x5_y13 (.clk(clknet_5_22__leaf_clk),
    .d(\state[197] ),
    .dl(\state[196] ),
    .dr(\state[198] ),
    .in_data(net12),
    .l(\state[212] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[213] ),
    .prev_out_data(\cell_outs[229] ),
    .r(\state[214] ),
    .reset(net77),
    .run(net60),
    .shift(net92),
    .state(\state[213] ),
    .u(\state[229] ),
    .ul(\state[228] ),
    .ur(\state[230] ));
 life_cell arr_cell_x5_y14 (.clk(clknet_5_23__leaf_clk),
    .d(\state[213] ),
    .dl(\state[212] ),
    .dr(\state[214] ),
    .in_data(net12),
    .l(\state[228] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[229] ),
    .prev_out_data(\cell_outs[245] ),
    .r(\state[230] ),
    .reset(net77),
    .run(net59),
    .shift(net92),
    .state(\state[229] ),
    .u(\state[245] ),
    .ul(\state[244] ),
    .ur(\state[246] ));
 life_cell arr_cell_x5_y15 (.clk(clknet_5_23__leaf_clk),
    .d(\state[229] ),
    .dl(\state[228] ),
    .dr(\state[230] ),
    .in_data(net12),
    .l(\state[244] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[245] ),
    .prev_out_data(net295),
    .r(\state[246] ),
    .reset(net77),
    .run(net58),
    .shift(net92),
    .state(\state[245] ),
    .u(net296),
    .ul(net297),
    .ur(net298));
 life_cell arr_cell_x5_y2 (.clk(clknet_5_3__leaf_clk),
    .d(\state[21] ),
    .dl(\state[20] ),
    .dr(\state[22] ),
    .in_data(net12),
    .l(\state[36] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[37] ),
    .prev_out_data(\cell_outs[53] ),
    .r(\state[38] ),
    .reset(net77),
    .run(net54),
    .shift(net92),
    .state(\state[37] ),
    .u(\state[53] ),
    .ul(\state[52] ),
    .ur(\state[54] ));
 life_cell arr_cell_x5_y3 (.clk(clknet_5_3__leaf_clk),
    .d(\state[37] ),
    .dl(\state[36] ),
    .dr(\state[38] ),
    .in_data(net12),
    .l(\state[52] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[53] ),
    .prev_out_data(\cell_outs[69] ),
    .r(\state[54] ),
    .reset(net77),
    .run(net55),
    .shift(net92),
    .state(\state[53] ),
    .u(\state[69] ),
    .ul(\state[68] ),
    .ur(\state[70] ));
 life_cell arr_cell_x5_y4 (.clk(clknet_5_6__leaf_clk),
    .d(\state[53] ),
    .dl(\state[52] ),
    .dr(\state[54] ),
    .in_data(net12),
    .l(\state[68] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[69] ),
    .prev_out_data(\cell_outs[85] ),
    .r(\state[70] ),
    .reset(net77),
    .run(net56),
    .shift(net92),
    .state(\state[69] ),
    .u(\state[85] ),
    .ul(\state[84] ),
    .ur(\state[86] ));
 life_cell arr_cell_x5_y5 (.clk(clknet_5_6__leaf_clk),
    .d(\state[69] ),
    .dl(\state[68] ),
    .dr(\state[70] ),
    .in_data(net12),
    .l(\state[84] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[85] ),
    .prev_out_data(\cell_outs[101] ),
    .r(\state[86] ),
    .reset(net77),
    .run(net57),
    .shift(net92),
    .state(\state[85] ),
    .u(\state[101] ),
    .ul(\state[100] ),
    .ur(\state[102] ));
 life_cell arr_cell_x5_y6 (.clk(clknet_5_7__leaf_clk),
    .d(\state[85] ),
    .dl(\state[84] ),
    .dr(\state[86] ),
    .in_data(net12),
    .l(\state[100] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[101] ),
    .prev_out_data(\cell_outs[117] ),
    .r(\state[102] ),
    .reset(net77),
    .run(net66),
    .shift(net92),
    .state(\state[101] ),
    .u(\state[117] ),
    .ul(\state[116] ),
    .ur(\state[118] ));
 life_cell arr_cell_x5_y7 (.clk(clknet_5_7__leaf_clk),
    .d(\state[101] ),
    .dl(\state[100] ),
    .dr(\state[102] ),
    .in_data(net12),
    .l(\state[116] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[117] ),
    .prev_out_data(\cell_outs[133] ),
    .r(\state[118] ),
    .reset(net77),
    .run(net25),
    .shift(net92),
    .state(\state[117] ),
    .u(\state[133] ),
    .ul(\state[132] ),
    .ur(\state[134] ));
 life_cell arr_cell_x5_y8 (.clk(clknet_5_18__leaf_clk),
    .d(\state[117] ),
    .dl(\state[116] ),
    .dr(\state[118] ),
    .in_data(net12),
    .l(\state[132] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[133] ),
    .prev_out_data(\cell_outs[149] ),
    .r(\state[134] ),
    .reset(net77),
    .run(net65),
    .shift(net92),
    .state(\state[133] ),
    .u(\state[149] ),
    .ul(\state[148] ),
    .ur(\state[150] ));
 life_cell arr_cell_x5_y9 (.clk(clknet_5_18__leaf_clk),
    .d(\state[133] ),
    .dl(\state[132] ),
    .dr(\state[134] ),
    .in_data(net12),
    .l(\state[148] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[149] ),
    .prev_out_data(\cell_outs[165] ),
    .r(\state[150] ),
    .reset(net77),
    .run(net64),
    .shift(net92),
    .state(\state[149] ),
    .u(\state[165] ),
    .ul(\state[164] ),
    .ur(\state[166] ));
 life_cell arr_cell_x6_y0 (.clk(clknet_5_2__leaf_clk),
    .d(net299),
    .dl(net300),
    .dr(net301),
    .in_data(net13),
    .l(\state[5] ),
    .load_in(net46),
    .load_out(net22),
    .out_data(\cell_outs[6] ),
    .prev_out_data(\cell_outs[22] ),
    .r(\state[7] ),
    .reset(net76),
    .run(net52),
    .shift(net91),
    .state(\state[6] ),
    .u(\state[22] ),
    .ul(\state[21] ),
    .ur(\state[23] ));
 life_cell arr_cell_x6_y1 (.clk(clknet_5_2__leaf_clk),
    .d(\state[6] ),
    .dl(\state[5] ),
    .dr(\state[7] ),
    .in_data(net13),
    .l(\state[21] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[22] ),
    .prev_out_data(\cell_outs[38] ),
    .r(\state[23] ),
    .reset(net76),
    .run(net53),
    .shift(net91),
    .state(\state[22] ),
    .u(\state[38] ),
    .ul(\state[37] ),
    .ur(\state[39] ));
 life_cell arr_cell_x6_y10 (.clk(clknet_5_19__leaf_clk),
    .d(\state[150] ),
    .dl(\state[149] ),
    .dr(\state[151] ),
    .in_data(net13),
    .l(\state[165] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[166] ),
    .prev_out_data(\cell_outs[182] ),
    .r(\state[167] ),
    .reset(net76),
    .run(net63),
    .shift(net91),
    .state(\state[166] ),
    .u(\state[182] ),
    .ul(\state[181] ),
    .ur(\state[183] ));
 life_cell arr_cell_x6_y11 (.clk(clknet_5_19__leaf_clk),
    .d(\state[166] ),
    .dl(\state[165] ),
    .dr(\state[167] ),
    .in_data(net13),
    .l(\state[181] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[182] ),
    .prev_out_data(\cell_outs[198] ),
    .r(\state[183] ),
    .reset(net76),
    .run(net62),
    .shift(net91),
    .state(\state[182] ),
    .u(\state[198] ),
    .ul(\state[197] ),
    .ur(\state[199] ));
 life_cell arr_cell_x6_y12 (.clk(clknet_5_22__leaf_clk),
    .d(\state[182] ),
    .dl(\state[181] ),
    .dr(\state[183] ),
    .in_data(net13),
    .l(\state[197] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[198] ),
    .prev_out_data(\cell_outs[214] ),
    .r(\state[199] ),
    .reset(net76),
    .run(net61),
    .shift(net91),
    .state(\state[198] ),
    .u(\state[214] ),
    .ul(\state[213] ),
    .ur(\state[215] ));
 life_cell arr_cell_x6_y13 (.clk(clknet_5_22__leaf_clk),
    .d(\state[198] ),
    .dl(\state[197] ),
    .dr(\state[199] ),
    .in_data(net13),
    .l(\state[213] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[214] ),
    .prev_out_data(\cell_outs[230] ),
    .r(\state[215] ),
    .reset(net76),
    .run(net60),
    .shift(net91),
    .state(\state[214] ),
    .u(\state[230] ),
    .ul(\state[229] ),
    .ur(\state[231] ));
 life_cell arr_cell_x6_y14 (.clk(clknet_5_23__leaf_clk),
    .d(\state[214] ),
    .dl(\state[213] ),
    .dr(\state[215] ),
    .in_data(net13),
    .l(\state[229] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[230] ),
    .prev_out_data(\cell_outs[246] ),
    .r(\state[231] ),
    .reset(net76),
    .run(net59),
    .shift(net91),
    .state(\state[230] ),
    .u(\state[246] ),
    .ul(\state[245] ),
    .ur(\state[247] ));
 life_cell arr_cell_x6_y15 (.clk(clknet_5_23__leaf_clk),
    .d(\state[230] ),
    .dl(\state[229] ),
    .dr(\state[231] ),
    .in_data(net13),
    .l(\state[245] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[246] ),
    .prev_out_data(net302),
    .r(\state[247] ),
    .reset(net76),
    .run(net58),
    .shift(net91),
    .state(\state[246] ),
    .u(net303),
    .ul(net304),
    .ur(net305));
 life_cell arr_cell_x6_y2 (.clk(clknet_5_3__leaf_clk),
    .d(\state[22] ),
    .dl(\state[21] ),
    .dr(\state[23] ),
    .in_data(net13),
    .l(\state[37] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[38] ),
    .prev_out_data(\cell_outs[54] ),
    .r(\state[39] ),
    .reset(net76),
    .run(net54),
    .shift(net91),
    .state(\state[38] ),
    .u(\state[54] ),
    .ul(\state[53] ),
    .ur(\state[55] ));
 life_cell arr_cell_x6_y3 (.clk(clknet_5_3__leaf_clk),
    .d(\state[38] ),
    .dl(\state[37] ),
    .dr(\state[39] ),
    .in_data(net13),
    .l(\state[53] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[54] ),
    .prev_out_data(\cell_outs[70] ),
    .r(\state[55] ),
    .reset(net76),
    .run(net55),
    .shift(net91),
    .state(\state[54] ),
    .u(\state[70] ),
    .ul(\state[69] ),
    .ur(\state[71] ));
 life_cell arr_cell_x6_y4 (.clk(clknet_5_6__leaf_clk),
    .d(\state[54] ),
    .dl(\state[53] ),
    .dr(\state[55] ),
    .in_data(net13),
    .l(\state[69] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[70] ),
    .prev_out_data(\cell_outs[86] ),
    .r(\state[71] ),
    .reset(net76),
    .run(net56),
    .shift(net91),
    .state(\state[70] ),
    .u(\state[86] ),
    .ul(\state[85] ),
    .ur(\state[87] ));
 life_cell arr_cell_x6_y5 (.clk(clknet_5_6__leaf_clk),
    .d(\state[70] ),
    .dl(\state[69] ),
    .dr(\state[71] ),
    .in_data(net13),
    .l(\state[85] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[86] ),
    .prev_out_data(\cell_outs[102] ),
    .r(\state[87] ),
    .reset(net76),
    .run(net57),
    .shift(net91),
    .state(\state[86] ),
    .u(\state[102] ),
    .ul(\state[101] ),
    .ur(\state[103] ));
 life_cell arr_cell_x6_y6 (.clk(clknet_5_7__leaf_clk),
    .d(\state[86] ),
    .dl(\state[85] ),
    .dr(\state[87] ),
    .in_data(net13),
    .l(\state[101] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[102] ),
    .prev_out_data(\cell_outs[118] ),
    .r(\state[103] ),
    .reset(net76),
    .run(net66),
    .shift(net91),
    .state(\state[102] ),
    .u(\state[118] ),
    .ul(\state[117] ),
    .ur(\state[119] ));
 life_cell arr_cell_x6_y7 (.clk(clknet_5_7__leaf_clk),
    .d(\state[102] ),
    .dl(\state[101] ),
    .dr(\state[103] ),
    .in_data(net13),
    .l(\state[117] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[118] ),
    .prev_out_data(\cell_outs[134] ),
    .r(\state[119] ),
    .reset(net76),
    .run(net25),
    .shift(net91),
    .state(\state[118] ),
    .u(\state[134] ),
    .ul(\state[133] ),
    .ur(\state[135] ));
 life_cell arr_cell_x6_y8 (.clk(clknet_5_18__leaf_clk),
    .d(\state[118] ),
    .dl(\state[117] ),
    .dr(\state[119] ),
    .in_data(net13),
    .l(\state[133] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[134] ),
    .prev_out_data(\cell_outs[150] ),
    .r(\state[135] ),
    .reset(net76),
    .run(net65),
    .shift(net91),
    .state(\state[134] ),
    .u(\state[150] ),
    .ul(\state[149] ),
    .ur(\state[151] ));
 life_cell arr_cell_x6_y9 (.clk(clknet_5_18__leaf_clk),
    .d(\state[134] ),
    .dl(\state[133] ),
    .dr(\state[135] ),
    .in_data(net13),
    .l(\state[149] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[150] ),
    .prev_out_data(\cell_outs[166] ),
    .r(\state[151] ),
    .reset(net76),
    .run(net64),
    .shift(net91),
    .state(\state[150] ),
    .u(\state[166] ),
    .ul(\state[165] ),
    .ur(\state[167] ));
 life_cell arr_cell_x7_y0 (.clk(clknet_5_2__leaf_clk),
    .d(net306),
    .dl(net307),
    .dr(net308),
    .in_data(net14),
    .l(\state[6] ),
    .load_in(net46),
    .load_out(net22),
    .out_data(\cell_outs[7] ),
    .prev_out_data(\cell_outs[23] ),
    .r(\state[8] ),
    .reset(net75),
    .run(net52),
    .shift(net90),
    .state(\state[7] ),
    .u(\state[23] ),
    .ul(\state[22] ),
    .ur(\state[24] ));
 life_cell arr_cell_x7_y1 (.clk(clknet_5_2__leaf_clk),
    .d(\state[7] ),
    .dl(\state[6] ),
    .dr(\state[8] ),
    .in_data(net14),
    .l(\state[22] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[23] ),
    .prev_out_data(\cell_outs[39] ),
    .r(\state[24] ),
    .reset(net75),
    .run(net53),
    .shift(net90),
    .state(\state[23] ),
    .u(\state[39] ),
    .ul(\state[38] ),
    .ur(\state[40] ));
 life_cell arr_cell_x7_y10 (.clk(clknet_5_19__leaf_clk),
    .d(\state[151] ),
    .dl(\state[150] ),
    .dr(\state[152] ),
    .in_data(net14),
    .l(\state[166] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[167] ),
    .prev_out_data(\cell_outs[183] ),
    .r(\state[168] ),
    .reset(net75),
    .run(net63),
    .shift(net90),
    .state(\state[167] ),
    .u(\state[183] ),
    .ul(\state[182] ),
    .ur(\state[184] ));
 life_cell arr_cell_x7_y11 (.clk(clknet_5_19__leaf_clk),
    .d(\state[167] ),
    .dl(\state[166] ),
    .dr(\state[168] ),
    .in_data(net14),
    .l(\state[182] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[183] ),
    .prev_out_data(\cell_outs[199] ),
    .r(\state[184] ),
    .reset(net75),
    .run(net62),
    .shift(net90),
    .state(\state[183] ),
    .u(\state[199] ),
    .ul(\state[198] ),
    .ur(\state[200] ));
 life_cell arr_cell_x7_y12 (.clk(clknet_5_22__leaf_clk),
    .d(\state[183] ),
    .dl(\state[182] ),
    .dr(\state[184] ),
    .in_data(net14),
    .l(\state[198] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[199] ),
    .prev_out_data(\cell_outs[215] ),
    .r(\state[200] ),
    .reset(net75),
    .run(net61),
    .shift(net90),
    .state(\state[199] ),
    .u(\state[215] ),
    .ul(\state[214] ),
    .ur(\state[216] ));
 life_cell arr_cell_x7_y13 (.clk(clknet_5_22__leaf_clk),
    .d(\state[199] ),
    .dl(\state[198] ),
    .dr(\state[200] ),
    .in_data(net14),
    .l(\state[214] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[215] ),
    .prev_out_data(\cell_outs[231] ),
    .r(\state[216] ),
    .reset(net75),
    .run(net60),
    .shift(net90),
    .state(\state[215] ),
    .u(\state[231] ),
    .ul(\state[230] ),
    .ur(\state[232] ));
 life_cell arr_cell_x7_y14 (.clk(clknet_5_23__leaf_clk),
    .d(\state[215] ),
    .dl(\state[214] ),
    .dr(\state[216] ),
    .in_data(net14),
    .l(\state[230] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[231] ),
    .prev_out_data(\cell_outs[247] ),
    .r(\state[232] ),
    .reset(net75),
    .run(net59),
    .shift(net90),
    .state(\state[231] ),
    .u(\state[247] ),
    .ul(\state[246] ),
    .ur(\state[248] ));
 life_cell arr_cell_x7_y15 (.clk(clknet_5_23__leaf_clk),
    .d(\state[231] ),
    .dl(\state[230] ),
    .dr(\state[232] ),
    .in_data(net14),
    .l(\state[246] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[247] ),
    .prev_out_data(net309),
    .r(\state[248] ),
    .reset(net75),
    .run(net58),
    .shift(net90),
    .state(\state[247] ),
    .u(net310),
    .ul(net311),
    .ur(net312));
 life_cell arr_cell_x7_y2 (.clk(clknet_5_3__leaf_clk),
    .d(\state[23] ),
    .dl(\state[22] ),
    .dr(\state[24] ),
    .in_data(net14),
    .l(\state[38] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[39] ),
    .prev_out_data(\cell_outs[55] ),
    .r(\state[40] ),
    .reset(net75),
    .run(net54),
    .shift(net90),
    .state(\state[39] ),
    .u(\state[55] ),
    .ul(\state[54] ),
    .ur(\state[56] ));
 life_cell arr_cell_x7_y3 (.clk(clknet_5_3__leaf_clk),
    .d(\state[39] ),
    .dl(\state[38] ),
    .dr(\state[40] ),
    .in_data(net14),
    .l(\state[54] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[55] ),
    .prev_out_data(\cell_outs[71] ),
    .r(\state[56] ),
    .reset(net75),
    .run(net55),
    .shift(net90),
    .state(\state[55] ),
    .u(\state[71] ),
    .ul(\state[70] ),
    .ur(\state[72] ));
 life_cell arr_cell_x7_y4 (.clk(clknet_5_6__leaf_clk),
    .d(\state[55] ),
    .dl(\state[54] ),
    .dr(\state[56] ),
    .in_data(net14),
    .l(\state[70] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[71] ),
    .prev_out_data(\cell_outs[87] ),
    .r(\state[72] ),
    .reset(net75),
    .run(net56),
    .shift(net90),
    .state(\state[71] ),
    .u(\state[87] ),
    .ul(\state[86] ),
    .ur(\state[88] ));
 life_cell arr_cell_x7_y5 (.clk(clknet_5_6__leaf_clk),
    .d(\state[71] ),
    .dl(\state[70] ),
    .dr(\state[72] ),
    .in_data(net14),
    .l(\state[86] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[87] ),
    .prev_out_data(\cell_outs[103] ),
    .r(\state[88] ),
    .reset(net75),
    .run(net57),
    .shift(net90),
    .state(\state[87] ),
    .u(\state[103] ),
    .ul(\state[102] ),
    .ur(\state[104] ));
 life_cell arr_cell_x7_y6 (.clk(clknet_5_7__leaf_clk),
    .d(\state[87] ),
    .dl(\state[86] ),
    .dr(\state[88] ),
    .in_data(net14),
    .l(\state[102] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[103] ),
    .prev_out_data(\cell_outs[119] ),
    .r(\state[104] ),
    .reset(net75),
    .run(net66),
    .shift(net90),
    .state(\state[103] ),
    .u(\state[119] ),
    .ul(\state[118] ),
    .ur(\state[120] ));
 life_cell arr_cell_x7_y7 (.clk(clknet_5_7__leaf_clk),
    .d(\state[103] ),
    .dl(\state[102] ),
    .dr(\state[104] ),
    .in_data(net14),
    .l(\state[118] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[119] ),
    .prev_out_data(\cell_outs[135] ),
    .r(\state[120] ),
    .reset(net75),
    .run(net25),
    .shift(net90),
    .state(\state[119] ),
    .u(\state[135] ),
    .ul(\state[134] ),
    .ur(\state[136] ));
 life_cell arr_cell_x7_y8 (.clk(clknet_5_18__leaf_clk),
    .d(\state[119] ),
    .dl(\state[118] ),
    .dr(\state[120] ),
    .in_data(net14),
    .l(\state[134] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[135] ),
    .prev_out_data(\cell_outs[151] ),
    .r(\state[136] ),
    .reset(net75),
    .run(net65),
    .shift(net90),
    .state(\state[135] ),
    .u(\state[151] ),
    .ul(\state[150] ),
    .ur(\state[152] ));
 life_cell arr_cell_x7_y9 (.clk(clknet_5_18__leaf_clk),
    .d(\state[135] ),
    .dl(\state[134] ),
    .dr(\state[136] ),
    .in_data(net14),
    .l(\state[150] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[151] ),
    .prev_out_data(\cell_outs[167] ),
    .r(\state[152] ),
    .reset(net75),
    .run(net64),
    .shift(net90),
    .state(\state[151] ),
    .u(\state[167] ),
    .ul(\state[166] ),
    .ur(\state[168] ));
 life_cell arr_cell_x8_y0 (.clk(clknet_5_8__leaf_clk),
    .d(net313),
    .dl(net314),
    .dr(net315),
    .in_data(net15),
    .l(\state[7] ),
    .load_in(net45),
    .load_out(net22),
    .out_data(\cell_outs[8] ),
    .prev_out_data(\cell_outs[24] ),
    .r(\state[9] ),
    .reset(net74),
    .run(net52),
    .shift(net89),
    .state(\state[8] ),
    .u(\state[24] ),
    .ul(\state[23] ),
    .ur(\state[25] ));
 life_cell arr_cell_x8_y1 (.clk(clknet_5_8__leaf_clk),
    .d(\state[8] ),
    .dl(\state[7] ),
    .dr(\state[9] ),
    .in_data(net15),
    .l(\state[23] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[24] ),
    .prev_out_data(\cell_outs[40] ),
    .r(\state[25] ),
    .reset(net74),
    .run(net53),
    .shift(net89),
    .state(\state[24] ),
    .u(\state[40] ),
    .ul(\state[39] ),
    .ur(\state[41] ));
 life_cell arr_cell_x8_y10 (.clk(clknet_5_25__leaf_clk),
    .d(\state[152] ),
    .dl(\state[151] ),
    .dr(\state[153] ),
    .in_data(net15),
    .l(\state[167] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[168] ),
    .prev_out_data(\cell_outs[184] ),
    .r(\state[169] ),
    .reset(net74),
    .run(net63),
    .shift(net89),
    .state(\state[168] ),
    .u(\state[184] ),
    .ul(\state[183] ),
    .ur(\state[185] ));
 life_cell arr_cell_x8_y11 (.clk(clknet_5_25__leaf_clk),
    .d(\state[168] ),
    .dl(\state[167] ),
    .dr(\state[169] ),
    .in_data(net15),
    .l(\state[183] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[184] ),
    .prev_out_data(\cell_outs[200] ),
    .r(\state[185] ),
    .reset(net74),
    .run(net62),
    .shift(net89),
    .state(\state[184] ),
    .u(\state[200] ),
    .ul(\state[199] ),
    .ur(\state[201] ));
 life_cell arr_cell_x8_y12 (.clk(clknet_5_28__leaf_clk),
    .d(\state[184] ),
    .dl(\state[183] ),
    .dr(\state[185] ),
    .in_data(net15),
    .l(\state[199] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[200] ),
    .prev_out_data(\cell_outs[216] ),
    .r(\state[201] ),
    .reset(net74),
    .run(net61),
    .shift(net89),
    .state(\state[200] ),
    .u(\state[216] ),
    .ul(\state[215] ),
    .ur(\state[217] ));
 life_cell arr_cell_x8_y13 (.clk(clknet_5_28__leaf_clk),
    .d(\state[200] ),
    .dl(\state[199] ),
    .dr(\state[201] ),
    .in_data(net15),
    .l(\state[215] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[216] ),
    .prev_out_data(\cell_outs[232] ),
    .r(\state[217] ),
    .reset(net74),
    .run(net60),
    .shift(net89),
    .state(\state[216] ),
    .u(\state[232] ),
    .ul(\state[231] ),
    .ur(\state[233] ));
 life_cell arr_cell_x8_y14 (.clk(clknet_5_29__leaf_clk),
    .d(\state[216] ),
    .dl(\state[215] ),
    .dr(\state[217] ),
    .in_data(net15),
    .l(\state[231] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[232] ),
    .prev_out_data(\cell_outs[248] ),
    .r(\state[233] ),
    .reset(net74),
    .run(net59),
    .shift(net89),
    .state(\state[232] ),
    .u(\state[248] ),
    .ul(\state[247] ),
    .ur(\state[249] ));
 life_cell arr_cell_x8_y15 (.clk(clknet_5_29__leaf_clk),
    .d(\state[232] ),
    .dl(\state[231] ),
    .dr(\state[233] ),
    .in_data(net15),
    .l(\state[247] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[248] ),
    .prev_out_data(net316),
    .r(\state[249] ),
    .reset(net74),
    .run(net58),
    .shift(net89),
    .state(\state[248] ),
    .u(net317),
    .ul(net318),
    .ur(net319));
 life_cell arr_cell_x8_y2 (.clk(clknet_5_9__leaf_clk),
    .d(\state[24] ),
    .dl(\state[23] ),
    .dr(\state[25] ),
    .in_data(net15),
    .l(\state[39] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[40] ),
    .prev_out_data(\cell_outs[56] ),
    .r(\state[41] ),
    .reset(net74),
    .run(net54),
    .shift(net89),
    .state(\state[40] ),
    .u(\state[56] ),
    .ul(\state[55] ),
    .ur(\state[57] ));
 life_cell arr_cell_x8_y3 (.clk(clknet_5_9__leaf_clk),
    .d(\state[40] ),
    .dl(\state[39] ),
    .dr(\state[41] ),
    .in_data(net15),
    .l(\state[55] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[56] ),
    .prev_out_data(\cell_outs[72] ),
    .r(\state[57] ),
    .reset(net74),
    .run(net55),
    .shift(net89),
    .state(\state[56] ),
    .u(\state[72] ),
    .ul(\state[71] ),
    .ur(\state[73] ));
 life_cell arr_cell_x8_y4 (.clk(clknet_5_12__leaf_clk),
    .d(\state[56] ),
    .dl(\state[55] ),
    .dr(\state[57] ),
    .in_data(net15),
    .l(\state[71] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[72] ),
    .prev_out_data(\cell_outs[88] ),
    .r(\state[73] ),
    .reset(net74),
    .run(net56),
    .shift(net89),
    .state(\state[72] ),
    .u(\state[88] ),
    .ul(\state[87] ),
    .ur(\state[89] ));
 life_cell arr_cell_x8_y5 (.clk(clknet_5_12__leaf_clk),
    .d(\state[72] ),
    .dl(\state[71] ),
    .dr(\state[73] ),
    .in_data(net15),
    .l(\state[87] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[88] ),
    .prev_out_data(\cell_outs[104] ),
    .r(\state[89] ),
    .reset(net74),
    .run(net57),
    .shift(net89),
    .state(\state[88] ),
    .u(\state[104] ),
    .ul(\state[103] ),
    .ur(\state[105] ));
 life_cell arr_cell_x8_y6 (.clk(clknet_5_13__leaf_clk),
    .d(\state[88] ),
    .dl(\state[87] ),
    .dr(\state[89] ),
    .in_data(net15),
    .l(\state[103] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[104] ),
    .prev_out_data(\cell_outs[120] ),
    .r(\state[105] ),
    .reset(net74),
    .run(net66),
    .shift(net89),
    .state(\state[104] ),
    .u(\state[120] ),
    .ul(\state[119] ),
    .ur(\state[121] ));
 life_cell arr_cell_x8_y7 (.clk(clknet_5_13__leaf_clk),
    .d(\state[104] ),
    .dl(\state[103] ),
    .dr(\state[105] ),
    .in_data(net15),
    .l(\state[119] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[120] ),
    .prev_out_data(\cell_outs[136] ),
    .r(\state[121] ),
    .reset(net74),
    .run(net25),
    .shift(net89),
    .state(\state[120] ),
    .u(\state[136] ),
    .ul(\state[135] ),
    .ur(\state[137] ));
 life_cell arr_cell_x8_y8 (.clk(clknet_5_24__leaf_clk),
    .d(\state[120] ),
    .dl(\state[119] ),
    .dr(\state[121] ),
    .in_data(net15),
    .l(\state[135] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[136] ),
    .prev_out_data(\cell_outs[152] ),
    .r(\state[137] ),
    .reset(net74),
    .run(net65),
    .shift(net89),
    .state(\state[136] ),
    .u(\state[152] ),
    .ul(\state[151] ),
    .ur(\state[153] ));
 life_cell arr_cell_x8_y9 (.clk(clknet_5_24__leaf_clk),
    .d(\state[136] ),
    .dl(\state[135] ),
    .dr(\state[137] ),
    .in_data(net15),
    .l(\state[151] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[152] ),
    .prev_out_data(\cell_outs[168] ),
    .r(\state[153] ),
    .reset(net74),
    .run(net64),
    .shift(net89),
    .state(\state[152] ),
    .u(\state[168] ),
    .ul(\state[167] ),
    .ur(\state[169] ));
 life_cell arr_cell_x9_y0 (.clk(clknet_5_8__leaf_clk),
    .d(net320),
    .dl(net321),
    .dr(net322),
    .in_data(net16),
    .l(\state[8] ),
    .load_in(net45),
    .load_out(net22),
    .out_data(\cell_outs[9] ),
    .prev_out_data(\cell_outs[25] ),
    .r(\state[10] ),
    .reset(net73),
    .run(net52),
    .shift(net88),
    .state(\state[9] ),
    .u(\state[25] ),
    .ul(\state[24] ),
    .ur(\state[26] ));
 life_cell arr_cell_x9_y1 (.clk(clknet_5_8__leaf_clk),
    .d(\state[9] ),
    .dl(\state[8] ),
    .dr(\state[10] ),
    .in_data(net16),
    .l(\state[24] ),
    .load_in(_11_),
    .load_out(net115),
    .out_data(\cell_outs[25] ),
    .prev_out_data(\cell_outs[41] ),
    .r(\state[26] ),
    .reset(net73),
    .run(net53),
    .shift(net88),
    .state(\state[25] ),
    .u(\state[41] ),
    .ul(\state[40] ),
    .ur(\state[42] ));
 life_cell arr_cell_x9_y10 (.clk(clknet_5_25__leaf_clk),
    .d(\state[153] ),
    .dl(\state[152] ),
    .dr(\state[154] ),
    .in_data(net16),
    .l(\state[168] ),
    .load_in(_09_),
    .load_out(net102),
    .out_data(\cell_outs[169] ),
    .prev_out_data(\cell_outs[185] ),
    .r(\state[170] ),
    .reset(net73),
    .run(net63),
    .shift(net88),
    .state(\state[169] ),
    .u(\state[185] ),
    .ul(\state[184] ),
    .ur(\state[186] ));
 life_cell arr_cell_x9_y11 (.clk(clknet_5_25__leaf_clk),
    .d(\state[169] ),
    .dl(\state[168] ),
    .dr(\state[170] ),
    .in_data(net16),
    .l(\state[184] ),
    .load_in(_10_),
    .load_out(net101),
    .out_data(\cell_outs[185] ),
    .prev_out_data(\cell_outs[201] ),
    .r(\state[186] ),
    .reset(net73),
    .run(net62),
    .shift(net88),
    .state(\state[185] ),
    .u(\state[201] ),
    .ul(\state[200] ),
    .ur(\state[202] ));
 life_cell arr_cell_x9_y12 (.clk(clknet_5_28__leaf_clk),
    .d(\state[185] ),
    .dl(\state[184] ),
    .dr(\state[186] ),
    .in_data(net16),
    .l(\state[200] ),
    .load_in(_12_),
    .load_out(net100),
    .out_data(\cell_outs[201] ),
    .prev_out_data(\cell_outs[217] ),
    .r(\state[202] ),
    .reset(net73),
    .run(net61),
    .shift(net88),
    .state(\state[201] ),
    .u(\state[217] ),
    .ul(\state[216] ),
    .ur(\state[218] ));
 life_cell arr_cell_x9_y13 (.clk(clknet_5_28__leaf_clk),
    .d(\state[201] ),
    .dl(\state[200] ),
    .dr(\state[202] ),
    .in_data(net16),
    .l(\state[216] ),
    .load_in(_13_),
    .load_out(net99),
    .out_data(\cell_outs[217] ),
    .prev_out_data(\cell_outs[233] ),
    .r(\state[218] ),
    .reset(net73),
    .run(net60),
    .shift(net88),
    .state(\state[217] ),
    .u(\state[233] ),
    .ul(\state[232] ),
    .ur(\state[234] ));
 life_cell arr_cell_x9_y14 (.clk(clknet_5_29__leaf_clk),
    .d(\state[217] ),
    .dl(\state[216] ),
    .dr(\state[218] ),
    .in_data(net16),
    .l(\state[232] ),
    .load_in(_14_),
    .load_out(net98),
    .out_data(\cell_outs[233] ),
    .prev_out_data(\cell_outs[249] ),
    .r(\state[234] ),
    .reset(net73),
    .run(net59),
    .shift(net88),
    .state(\state[233] ),
    .u(\state[249] ),
    .ul(\state[248] ),
    .ur(\state[250] ));
 life_cell arr_cell_x9_y15 (.clk(clknet_5_29__leaf_clk),
    .d(\state[233] ),
    .dl(\state[232] ),
    .dr(\state[234] ),
    .in_data(net16),
    .l(\state[248] ),
    .load_in(_15_),
    .load_out(net97),
    .out_data(\cell_outs[249] ),
    .prev_out_data(net323),
    .r(\state[250] ),
    .reset(net73),
    .run(net58),
    .shift(net88),
    .state(\state[249] ),
    .u(net324),
    .ul(net325),
    .ur(net326));
 life_cell arr_cell_x9_y2 (.clk(clknet_5_9__leaf_clk),
    .d(\state[25] ),
    .dl(\state[24] ),
    .dr(\state[26] ),
    .in_data(net16),
    .l(\state[40] ),
    .load_in(_00_),
    .load_out(net110),
    .out_data(\cell_outs[41] ),
    .prev_out_data(\cell_outs[57] ),
    .r(\state[42] ),
    .reset(net73),
    .run(net54),
    .shift(net88),
    .state(\state[41] ),
    .u(\state[57] ),
    .ul(\state[56] ),
    .ur(\state[58] ));
 life_cell arr_cell_x9_y3 (.clk(clknet_5_9__leaf_clk),
    .d(\state[41] ),
    .dl(\state[40] ),
    .dr(\state[42] ),
    .in_data(net16),
    .l(\state[56] ),
    .load_in(_02_),
    .load_out(net109),
    .out_data(\cell_outs[57] ),
    .prev_out_data(\cell_outs[73] ),
    .r(\state[58] ),
    .reset(net73),
    .run(net55),
    .shift(net88),
    .state(\state[57] ),
    .u(\state[73] ),
    .ul(\state[72] ),
    .ur(\state[74] ));
 life_cell arr_cell_x9_y4 (.clk(clknet_5_12__leaf_clk),
    .d(\state[57] ),
    .dl(\state[56] ),
    .dr(\state[58] ),
    .in_data(net16),
    .l(\state[72] ),
    .load_in(_03_),
    .load_out(net108),
    .out_data(\cell_outs[73] ),
    .prev_out_data(\cell_outs[89] ),
    .r(\state[74] ),
    .reset(net73),
    .run(net56),
    .shift(net88),
    .state(\state[73] ),
    .u(\state[89] ),
    .ul(\state[88] ),
    .ur(\state[90] ));
 life_cell arr_cell_x9_y5 (.clk(clknet_5_12__leaf_clk),
    .d(\state[73] ),
    .dl(\state[72] ),
    .dr(\state[74] ),
    .in_data(net16),
    .l(\state[88] ),
    .load_in(_04_),
    .load_out(net107),
    .out_data(\cell_outs[89] ),
    .prev_out_data(\cell_outs[105] ),
    .r(\state[90] ),
    .reset(net73),
    .run(net57),
    .shift(net88),
    .state(\state[89] ),
    .u(\state[105] ),
    .ul(\state[104] ),
    .ur(\state[106] ));
 life_cell arr_cell_x9_y6 (.clk(clknet_5_13__leaf_clk),
    .d(\state[89] ),
    .dl(\state[88] ),
    .dr(\state[90] ),
    .in_data(net16),
    .l(\state[104] ),
    .load_in(_05_),
    .load_out(net106),
    .out_data(\cell_outs[105] ),
    .prev_out_data(\cell_outs[121] ),
    .r(\state[106] ),
    .reset(net73),
    .run(net66),
    .shift(net88),
    .state(\state[105] ),
    .u(\state[121] ),
    .ul(\state[120] ),
    .ur(\state[122] ));
 life_cell arr_cell_x9_y7 (.clk(clknet_5_13__leaf_clk),
    .d(\state[105] ),
    .dl(\state[104] ),
    .dr(\state[106] ),
    .in_data(net16),
    .l(\state[120] ),
    .load_in(_06_),
    .load_out(net105),
    .out_data(\cell_outs[121] ),
    .prev_out_data(\cell_outs[137] ),
    .r(\state[122] ),
    .reset(net73),
    .run(net25),
    .shift(net88),
    .state(\state[121] ),
    .u(\state[137] ),
    .ul(\state[136] ),
    .ur(\state[138] ));
 life_cell arr_cell_x9_y8 (.clk(clknet_5_24__leaf_clk),
    .d(\state[121] ),
    .dl(\state[120] ),
    .dr(\state[122] ),
    .in_data(net16),
    .l(\state[136] ),
    .load_in(_07_),
    .load_out(net104),
    .out_data(\cell_outs[137] ),
    .prev_out_data(\cell_outs[153] ),
    .r(\state[138] ),
    .reset(net73),
    .run(net65),
    .shift(net88),
    .state(\state[137] ),
    .u(\state[153] ),
    .ul(\state[152] ),
    .ur(\state[154] ));
 life_cell arr_cell_x9_y9 (.clk(clknet_5_24__leaf_clk),
    .d(\state[137] ),
    .dl(\state[136] ),
    .dr(\state[138] ),
    .in_data(net16),
    .l(\state[152] ),
    .load_in(_08_),
    .load_out(net103),
    .out_data(\cell_outs[153] ),
    .prev_out_data(\cell_outs[169] ),
    .r(\state[154] ),
    .reset(net73),
    .run(net64),
    .shift(net88),
    .state(\state[153] ),
    .u(\state[169] ),
    .ul(\state[168] ),
    .ur(\state[170] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__decap_3 PHY_1064 ();
 sky130_fd_sc_hd__decap_3 PHY_1065 ();
 sky130_fd_sc_hd__decap_3 PHY_1066 ();
 sky130_fd_sc_hd__decap_3 PHY_1067 ();
 sky130_fd_sc_hd__decap_3 PHY_1068 ();
 sky130_fd_sc_hd__decap_3 PHY_1069 ();
 sky130_fd_sc_hd__decap_3 PHY_1070 ();
 sky130_fd_sc_hd__decap_3 PHY_1071 ();
 sky130_fd_sc_hd__decap_3 PHY_1072 ();
 sky130_fd_sc_hd__decap_3 PHY_1073 ();
 sky130_fd_sc_hd__decap_3 PHY_1074 ();
 sky130_fd_sc_hd__decap_3 PHY_1075 ();
 sky130_fd_sc_hd__decap_3 PHY_1076 ();
 sky130_fd_sc_hd__decap_3 PHY_1077 ();
 sky130_fd_sc_hd__decap_3 PHY_1078 ();
 sky130_fd_sc_hd__decap_3 PHY_1079 ();
 sky130_fd_sc_hd__decap_3 PHY_1080 ();
 sky130_fd_sc_hd__decap_3 PHY_1081 ();
 sky130_fd_sc_hd__decap_3 PHY_1082 ();
 sky130_fd_sc_hd__decap_3 PHY_1083 ();
 sky130_fd_sc_hd__decap_3 PHY_1084 ();
 sky130_fd_sc_hd__decap_3 PHY_1085 ();
 sky130_fd_sc_hd__decap_3 PHY_1086 ();
 sky130_fd_sc_hd__decap_3 PHY_1087 ();
 sky130_fd_sc_hd__decap_3 PHY_1088 ();
 sky130_fd_sc_hd__decap_3 PHY_1089 ();
 sky130_fd_sc_hd__decap_3 PHY_1090 ();
 sky130_fd_sc_hd__decap_3 PHY_1091 ();
 sky130_fd_sc_hd__decap_3 PHY_1092 ();
 sky130_fd_sc_hd__decap_3 PHY_1093 ();
 sky130_fd_sc_hd__decap_3 PHY_1094 ();
 sky130_fd_sc_hd__decap_3 PHY_1095 ();
 sky130_fd_sc_hd__decap_3 PHY_1096 ();
 sky130_fd_sc_hd__decap_3 PHY_1097 ();
 sky130_fd_sc_hd__decap_3 PHY_1098 ();
 sky130_fd_sc_hd__decap_3 PHY_1099 ();
 sky130_fd_sc_hd__decap_3 PHY_1100 ();
 sky130_fd_sc_hd__decap_3 PHY_1101 ();
 sky130_fd_sc_hd__decap_3 PHY_1102 ();
 sky130_fd_sc_hd__decap_3 PHY_1103 ();
 sky130_fd_sc_hd__decap_3 PHY_1104 ();
 sky130_fd_sc_hd__decap_3 PHY_1105 ();
 sky130_fd_sc_hd__decap_3 PHY_1106 ();
 sky130_fd_sc_hd__decap_3 PHY_1107 ();
 sky130_fd_sc_hd__decap_3 PHY_1108 ();
 sky130_fd_sc_hd__decap_3 PHY_1109 ();
 sky130_fd_sc_hd__decap_3 PHY_1110 ();
 sky130_fd_sc_hd__decap_3 PHY_1111 ();
 sky130_fd_sc_hd__decap_3 PHY_1112 ();
 sky130_fd_sc_hd__decap_3 PHY_1113 ();
 sky130_fd_sc_hd__decap_3 PHY_1114 ();
 sky130_fd_sc_hd__decap_3 PHY_1115 ();
 sky130_fd_sc_hd__decap_3 PHY_1116 ();
 sky130_fd_sc_hd__decap_3 PHY_1117 ();
 sky130_fd_sc_hd__decap_3 PHY_1118 ();
 sky130_fd_sc_hd__decap_3 PHY_1119 ();
 sky130_fd_sc_hd__decap_3 PHY_1120 ();
 sky130_fd_sc_hd__decap_3 PHY_1121 ();
 sky130_fd_sc_hd__decap_3 PHY_1122 ();
 sky130_fd_sc_hd__decap_3 PHY_1123 ();
 sky130_fd_sc_hd__decap_3 PHY_1124 ();
 sky130_fd_sc_hd__decap_3 PHY_1125 ();
 sky130_fd_sc_hd__decap_3 PHY_1126 ();
 sky130_fd_sc_hd__decap_3 PHY_1127 ();
 sky130_fd_sc_hd__decap_3 PHY_1128 ();
 sky130_fd_sc_hd__decap_3 PHY_1129 ();
 sky130_fd_sc_hd__decap_3 PHY_1130 ();
 sky130_fd_sc_hd__decap_3 PHY_1131 ();
 sky130_fd_sc_hd__decap_3 PHY_1132 ();
 sky130_fd_sc_hd__decap_3 PHY_1133 ();
 sky130_fd_sc_hd__decap_3 PHY_1134 ();
 sky130_fd_sc_hd__decap_3 PHY_1135 ();
 sky130_fd_sc_hd__decap_3 PHY_1136 ();
 sky130_fd_sc_hd__decap_3 PHY_1137 ();
 sky130_fd_sc_hd__decap_3 PHY_1138 ();
 sky130_fd_sc_hd__decap_3 PHY_1139 ();
 sky130_fd_sc_hd__decap_3 PHY_1140 ();
 sky130_fd_sc_hd__decap_3 PHY_1141 ();
 sky130_fd_sc_hd__decap_3 PHY_1142 ();
 sky130_fd_sc_hd__decap_3 PHY_1143 ();
 sky130_fd_sc_hd__decap_3 PHY_1144 ();
 sky130_fd_sc_hd__decap_3 PHY_1145 ();
 sky130_fd_sc_hd__decap_3 PHY_1146 ();
 sky130_fd_sc_hd__decap_3 PHY_1147 ();
 sky130_fd_sc_hd__decap_3 PHY_1148 ();
 sky130_fd_sc_hd__decap_3 PHY_1149 ();
 sky130_fd_sc_hd__decap_3 PHY_1150 ();
 sky130_fd_sc_hd__decap_3 PHY_1151 ();
 sky130_fd_sc_hd__decap_3 PHY_1152 ();
 sky130_fd_sc_hd__decap_3 PHY_1153 ();
 sky130_fd_sc_hd__decap_3 PHY_1154 ();
 sky130_fd_sc_hd__decap_3 PHY_1155 ();
 sky130_fd_sc_hd__decap_3 PHY_1156 ();
 sky130_fd_sc_hd__decap_3 PHY_1157 ();
 sky130_fd_sc_hd__decap_3 PHY_1158 ();
 sky130_fd_sc_hd__decap_3 PHY_1159 ();
 sky130_fd_sc_hd__decap_3 PHY_1160 ();
 sky130_fd_sc_hd__decap_3 PHY_1161 ();
 sky130_fd_sc_hd__decap_3 PHY_1162 ();
 sky130_fd_sc_hd__decap_3 PHY_1163 ();
 sky130_fd_sc_hd__decap_3 PHY_1164 ();
 sky130_fd_sc_hd__decap_3 PHY_1165 ();
 sky130_fd_sc_hd__decap_3 PHY_1166 ();
 sky130_fd_sc_hd__decap_3 PHY_1167 ();
 sky130_fd_sc_hd__decap_3 PHY_1168 ();
 sky130_fd_sc_hd__decap_3 PHY_1169 ();
 sky130_fd_sc_hd__decap_3 PHY_1170 ();
 sky130_fd_sc_hd__decap_3 PHY_1171 ();
 sky130_fd_sc_hd__decap_3 PHY_1172 ();
 sky130_fd_sc_hd__decap_3 PHY_1173 ();
 sky130_fd_sc_hd__decap_3 PHY_1174 ();
 sky130_fd_sc_hd__decap_3 PHY_1175 ();
 sky130_fd_sc_hd__decap_3 PHY_1176 ();
 sky130_fd_sc_hd__decap_3 PHY_1177 ();
 sky130_fd_sc_hd__decap_3 PHY_1178 ();
 sky130_fd_sc_hd__decap_3 PHY_1179 ();
 sky130_fd_sc_hd__decap_3 PHY_1180 ();
 sky130_fd_sc_hd__decap_3 PHY_1181 ();
 sky130_fd_sc_hd__decap_3 PHY_1182 ();
 sky130_fd_sc_hd__decap_3 PHY_1183 ();
 sky130_fd_sc_hd__decap_3 PHY_1184 ();
 sky130_fd_sc_hd__decap_3 PHY_1185 ();
 sky130_fd_sc_hd__decap_3 PHY_1186 ();
 sky130_fd_sc_hd__decap_3 PHY_1187 ();
 sky130_fd_sc_hd__decap_3 PHY_1188 ();
 sky130_fd_sc_hd__decap_3 PHY_1189 ();
 sky130_fd_sc_hd__decap_3 PHY_1190 ();
 sky130_fd_sc_hd__decap_3 PHY_1191 ();
 sky130_fd_sc_hd__decap_3 PHY_1192 ();
 sky130_fd_sc_hd__decap_3 PHY_1193 ();
 sky130_fd_sc_hd__decap_3 PHY_1194 ();
 sky130_fd_sc_hd__decap_3 PHY_1195 ();
 sky130_fd_sc_hd__decap_3 PHY_1196 ();
 sky130_fd_sc_hd__decap_3 PHY_1197 ();
 sky130_fd_sc_hd__decap_3 PHY_1198 ();
 sky130_fd_sc_hd__decap_3 PHY_1199 ();
 sky130_fd_sc_hd__decap_3 PHY_1200 ();
 sky130_fd_sc_hd__decap_3 PHY_1201 ();
 sky130_fd_sc_hd__decap_3 PHY_1202 ();
 sky130_fd_sc_hd__decap_3 PHY_1203 ();
 sky130_fd_sc_hd__decap_3 PHY_1204 ();
 sky130_fd_sc_hd__decap_3 PHY_1205 ();
 sky130_fd_sc_hd__decap_3 PHY_1206 ();
 sky130_fd_sc_hd__decap_3 PHY_1207 ();
 sky130_fd_sc_hd__decap_3 PHY_1208 ();
 sky130_fd_sc_hd__decap_3 PHY_1209 ();
 sky130_fd_sc_hd__decap_3 PHY_1210 ();
 sky130_fd_sc_hd__decap_3 PHY_1211 ();
 sky130_fd_sc_hd__decap_3 PHY_1212 ();
 sky130_fd_sc_hd__decap_3 PHY_1213 ();
 sky130_fd_sc_hd__decap_3 PHY_1214 ();
 sky130_fd_sc_hd__decap_3 PHY_1215 ();
 sky130_fd_sc_hd__decap_3 PHY_1216 ();
 sky130_fd_sc_hd__decap_3 PHY_1217 ();
 sky130_fd_sc_hd__decap_3 PHY_1218 ();
 sky130_fd_sc_hd__decap_3 PHY_1219 ();
 sky130_fd_sc_hd__decap_3 PHY_1220 ();
 sky130_fd_sc_hd__decap_3 PHY_1221 ();
 sky130_fd_sc_hd__decap_3 PHY_1222 ();
 sky130_fd_sc_hd__decap_3 PHY_1223 ();
 sky130_fd_sc_hd__decap_3 PHY_1224 ();
 sky130_fd_sc_hd__decap_3 PHY_1225 ();
 sky130_fd_sc_hd__decap_3 PHY_1226 ();
 sky130_fd_sc_hd__decap_3 PHY_1227 ();
 sky130_fd_sc_hd__decap_3 PHY_1228 ();
 sky130_fd_sc_hd__decap_3 PHY_1229 ();
 sky130_fd_sc_hd__decap_3 PHY_1230 ();
 sky130_fd_sc_hd__decap_3 PHY_1231 ();
 sky130_fd_sc_hd__decap_3 PHY_1232 ();
 sky130_fd_sc_hd__decap_3 PHY_1233 ();
 sky130_fd_sc_hd__decap_3 PHY_1234 ();
 sky130_fd_sc_hd__decap_3 PHY_1235 ();
 sky130_fd_sc_hd__decap_3 PHY_1236 ();
 sky130_fd_sc_hd__decap_3 PHY_1237 ();
 sky130_fd_sc_hd__decap_3 PHY_1238 ();
 sky130_fd_sc_hd__decap_3 PHY_1239 ();
 sky130_fd_sc_hd__decap_3 PHY_1240 ();
 sky130_fd_sc_hd__decap_3 PHY_1241 ();
 sky130_fd_sc_hd__decap_3 PHY_1242 ();
 sky130_fd_sc_hd__decap_3 PHY_1243 ();
 sky130_fd_sc_hd__decap_3 PHY_1244 ();
 sky130_fd_sc_hd__decap_3 PHY_1245 ();
 sky130_fd_sc_hd__decap_3 PHY_1246 ();
 sky130_fd_sc_hd__decap_3 PHY_1247 ();
 sky130_fd_sc_hd__decap_3 PHY_1248 ();
 sky130_fd_sc_hd__decap_3 PHY_1249 ();
 sky130_fd_sc_hd__decap_3 PHY_1250 ();
 sky130_fd_sc_hd__decap_3 PHY_1251 ();
 sky130_fd_sc_hd__decap_3 PHY_1252 ();
 sky130_fd_sc_hd__decap_3 PHY_1253 ();
 sky130_fd_sc_hd__decap_3 PHY_1254 ();
 sky130_fd_sc_hd__decap_3 PHY_1255 ();
 sky130_fd_sc_hd__decap_3 PHY_1256 ();
 sky130_fd_sc_hd__decap_3 PHY_1257 ();
 sky130_fd_sc_hd__decap_3 PHY_1258 ();
 sky130_fd_sc_hd__decap_3 PHY_1259 ();
 sky130_fd_sc_hd__decap_3 PHY_1260 ();
 sky130_fd_sc_hd__decap_3 PHY_1261 ();
 sky130_fd_sc_hd__decap_3 PHY_1262 ();
 sky130_fd_sc_hd__decap_3 PHY_1263 ();
 sky130_fd_sc_hd__decap_3 PHY_1264 ();
 sky130_fd_sc_hd__decap_3 PHY_1265 ();
 sky130_fd_sc_hd__decap_3 PHY_1266 ();
 sky130_fd_sc_hd__decap_3 PHY_1267 ();
 sky130_fd_sc_hd__decap_3 PHY_1268 ();
 sky130_fd_sc_hd__decap_3 PHY_1269 ();
 sky130_fd_sc_hd__decap_3 PHY_1270 ();
 sky130_fd_sc_hd__decap_3 PHY_1271 ();
 sky130_fd_sc_hd__decap_3 PHY_1272 ();
 sky130_fd_sc_hd__decap_3 PHY_1273 ();
 sky130_fd_sc_hd__decap_3 PHY_1274 ();
 sky130_fd_sc_hd__decap_3 PHY_1275 ();
 sky130_fd_sc_hd__decap_3 PHY_1276 ();
 sky130_fd_sc_hd__decap_3 PHY_1277 ();
 sky130_fd_sc_hd__decap_3 PHY_1278 ();
 sky130_fd_sc_hd__decap_3 PHY_1279 ();
 sky130_fd_sc_hd__decap_3 PHY_1280 ();
 sky130_fd_sc_hd__decap_3 PHY_1281 ();
 sky130_fd_sc_hd__decap_3 PHY_1282 ();
 sky130_fd_sc_hd__decap_3 PHY_1283 ();
 sky130_fd_sc_hd__decap_3 PHY_1284 ();
 sky130_fd_sc_hd__decap_3 PHY_1285 ();
 sky130_fd_sc_hd__decap_3 PHY_1286 ();
 sky130_fd_sc_hd__decap_3 PHY_1287 ();
 sky130_fd_sc_hd__decap_3 PHY_1288 ();
 sky130_fd_sc_hd__decap_3 PHY_1289 ();
 sky130_fd_sc_hd__decap_3 PHY_1290 ();
 sky130_fd_sc_hd__decap_3 PHY_1291 ();
 sky130_fd_sc_hd__decap_3 PHY_1292 ();
 sky130_fd_sc_hd__decap_3 PHY_1293 ();
 sky130_fd_sc_hd__decap_3 PHY_1294 ();
 sky130_fd_sc_hd__decap_3 PHY_1295 ();
 sky130_fd_sc_hd__decap_3 PHY_1296 ();
 sky130_fd_sc_hd__decap_3 PHY_1297 ();
 sky130_fd_sc_hd__decap_3 PHY_1298 ();
 sky130_fd_sc_hd__decap_3 PHY_1299 ();
 sky130_fd_sc_hd__decap_3 PHY_1300 ();
 sky130_fd_sc_hd__decap_3 PHY_1301 ();
 sky130_fd_sc_hd__decap_3 PHY_1302 ();
 sky130_fd_sc_hd__decap_3 PHY_1303 ();
 sky130_fd_sc_hd__decap_3 PHY_1304 ();
 sky130_fd_sc_hd__decap_3 PHY_1305 ();
 sky130_fd_sc_hd__decap_3 PHY_1306 ();
 sky130_fd_sc_hd__decap_3 PHY_1307 ();
 sky130_fd_sc_hd__decap_3 PHY_1308 ();
 sky130_fd_sc_hd__decap_3 PHY_1309 ();
 sky130_fd_sc_hd__decap_3 PHY_1310 ();
 sky130_fd_sc_hd__decap_3 PHY_1311 ();
 sky130_fd_sc_hd__decap_3 PHY_1312 ();
 sky130_fd_sc_hd__decap_3 PHY_1313 ();
 sky130_fd_sc_hd__decap_3 PHY_1314 ();
 sky130_fd_sc_hd__decap_3 PHY_1315 ();
 sky130_fd_sc_hd__decap_3 PHY_1316 ();
 sky130_fd_sc_hd__decap_3 PHY_1317 ();
 sky130_fd_sc_hd__decap_3 PHY_1318 ();
 sky130_fd_sc_hd__decap_3 PHY_1319 ();
 sky130_fd_sc_hd__decap_3 PHY_1320 ();
 sky130_fd_sc_hd__decap_3 PHY_1321 ();
 sky130_fd_sc_hd__decap_3 PHY_1322 ();
 sky130_fd_sc_hd__decap_3 PHY_1323 ();
 sky130_fd_sc_hd__decap_3 PHY_1324 ();
 sky130_fd_sc_hd__decap_3 PHY_1325 ();
 sky130_fd_sc_hd__decap_3 PHY_1326 ();
 sky130_fd_sc_hd__decap_3 PHY_1327 ();
 sky130_fd_sc_hd__decap_3 PHY_1328 ();
 sky130_fd_sc_hd__decap_3 PHY_1329 ();
 sky130_fd_sc_hd__decap_3 PHY_1330 ();
 sky130_fd_sc_hd__decap_3 PHY_1331 ();
 sky130_fd_sc_hd__decap_3 PHY_1332 ();
 sky130_fd_sc_hd__decap_3 PHY_1333 ();
 sky130_fd_sc_hd__decap_3 PHY_1334 ();
 sky130_fd_sc_hd__decap_3 PHY_1335 ();
 sky130_fd_sc_hd__decap_3 PHY_1336 ();
 sky130_fd_sc_hd__decap_3 PHY_1337 ();
 sky130_fd_sc_hd__decap_3 PHY_1338 ();
 sky130_fd_sc_hd__decap_3 PHY_1339 ();
 sky130_fd_sc_hd__decap_3 PHY_1340 ();
 sky130_fd_sc_hd__decap_3 PHY_1341 ();
 sky130_fd_sc_hd__decap_3 PHY_1342 ();
 sky130_fd_sc_hd__decap_3 PHY_1343 ();
 sky130_fd_sc_hd__decap_3 PHY_1344 ();
 sky130_fd_sc_hd__decap_3 PHY_1345 ();
 sky130_fd_sc_hd__decap_3 PHY_1346 ();
 sky130_fd_sc_hd__decap_3 PHY_1347 ();
 sky130_fd_sc_hd__decap_3 PHY_1348 ();
 sky130_fd_sc_hd__decap_3 PHY_1349 ();
 sky130_fd_sc_hd__decap_3 PHY_1350 ();
 sky130_fd_sc_hd__decap_3 PHY_1351 ();
 sky130_fd_sc_hd__decap_3 PHY_1352 ();
 sky130_fd_sc_hd__decap_3 PHY_1353 ();
 sky130_fd_sc_hd__decap_3 PHY_1354 ();
 sky130_fd_sc_hd__decap_3 PHY_1355 ();
 sky130_fd_sc_hd__decap_3 PHY_1356 ();
 sky130_fd_sc_hd__decap_3 PHY_1357 ();
 sky130_fd_sc_hd__decap_3 PHY_1358 ();
 sky130_fd_sc_hd__decap_3 PHY_1359 ();
 sky130_fd_sc_hd__decap_3 PHY_1360 ();
 sky130_fd_sc_hd__decap_3 PHY_1361 ();
 sky130_fd_sc_hd__decap_3 PHY_1362 ();
 sky130_fd_sc_hd__decap_3 PHY_1363 ();
 sky130_fd_sc_hd__decap_3 PHY_1364 ();
 sky130_fd_sc_hd__decap_3 PHY_1365 ();
 sky130_fd_sc_hd__decap_3 PHY_1366 ();
 sky130_fd_sc_hd__decap_3 PHY_1367 ();
 sky130_fd_sc_hd__decap_3 PHY_1368 ();
 sky130_fd_sc_hd__decap_3 PHY_1369 ();
 sky130_fd_sc_hd__decap_3 PHY_1370 ();
 sky130_fd_sc_hd__decap_3 PHY_1371 ();
 sky130_fd_sc_hd__decap_3 PHY_1372 ();
 sky130_fd_sc_hd__decap_3 PHY_1373 ();
 sky130_fd_sc_hd__decap_3 PHY_1374 ();
 sky130_fd_sc_hd__decap_3 PHY_1375 ();
 sky130_fd_sc_hd__decap_3 PHY_1376 ();
 sky130_fd_sc_hd__decap_3 PHY_1377 ();
 sky130_fd_sc_hd__decap_3 PHY_1378 ();
 sky130_fd_sc_hd__decap_3 PHY_1379 ();
 sky130_fd_sc_hd__decap_3 PHY_1380 ();
 sky130_fd_sc_hd__decap_3 PHY_1381 ();
 sky130_fd_sc_hd__decap_3 PHY_1382 ();
 sky130_fd_sc_hd__decap_3 PHY_1383 ();
 sky130_fd_sc_hd__decap_3 PHY_1384 ();
 sky130_fd_sc_hd__decap_3 PHY_1385 ();
 sky130_fd_sc_hd__decap_3 PHY_1386 ();
 sky130_fd_sc_hd__decap_3 PHY_1387 ();
 sky130_fd_sc_hd__decap_3 PHY_1388 ();
 sky130_fd_sc_hd__decap_3 PHY_1389 ();
 sky130_fd_sc_hd__decap_3 PHY_1390 ();
 sky130_fd_sc_hd__decap_3 PHY_1391 ();
 sky130_fd_sc_hd__decap_3 PHY_1392 ();
 sky130_fd_sc_hd__decap_3 PHY_1393 ();
 sky130_fd_sc_hd__decap_3 PHY_1394 ();
 sky130_fd_sc_hd__decap_3 PHY_1395 ();
 sky130_fd_sc_hd__decap_3 PHY_1396 ();
 sky130_fd_sc_hd__decap_3 PHY_1397 ();
 sky130_fd_sc_hd__decap_3 PHY_1398 ();
 sky130_fd_sc_hd__decap_3 PHY_1399 ();
 sky130_fd_sc_hd__decap_3 PHY_1400 ();
 sky130_fd_sc_hd__decap_3 PHY_1401 ();
 sky130_fd_sc_hd__decap_3 PHY_1402 ();
 sky130_fd_sc_hd__decap_3 PHY_1403 ();
 sky130_fd_sc_hd__decap_3 PHY_1404 ();
 sky130_fd_sc_hd__decap_3 PHY_1405 ();
 sky130_fd_sc_hd__decap_3 PHY_1406 ();
 sky130_fd_sc_hd__decap_3 PHY_1407 ();
 sky130_fd_sc_hd__decap_3 PHY_1408 ();
 sky130_fd_sc_hd__decap_3 PHY_1409 ();
 sky130_fd_sc_hd__decap_3 PHY_1410 ();
 sky130_fd_sc_hd__decap_3 PHY_1411 ();
 sky130_fd_sc_hd__decap_3 PHY_1412 ();
 sky130_fd_sc_hd__decap_3 PHY_1413 ();
 sky130_fd_sc_hd__decap_3 PHY_1414 ();
 sky130_fd_sc_hd__decap_3 PHY_1415 ();
 sky130_fd_sc_hd__decap_3 PHY_1416 ();
 sky130_fd_sc_hd__decap_3 PHY_1417 ();
 sky130_fd_sc_hd__decap_3 PHY_1418 ();
 sky130_fd_sc_hd__decap_3 PHY_1419 ();
 sky130_fd_sc_hd__decap_3 PHY_1420 ();
 sky130_fd_sc_hd__decap_3 PHY_1421 ();
 sky130_fd_sc_hd__decap_3 PHY_1422 ();
 sky130_fd_sc_hd__decap_3 PHY_1423 ();
 sky130_fd_sc_hd__decap_3 PHY_1424 ();
 sky130_fd_sc_hd__decap_3 PHY_1425 ();
 sky130_fd_sc_hd__decap_3 PHY_1426 ();
 sky130_fd_sc_hd__decap_3 PHY_1427 ();
 sky130_fd_sc_hd__decap_3 PHY_1428 ();
 sky130_fd_sc_hd__decap_3 PHY_1429 ();
 sky130_fd_sc_hd__decap_3 PHY_1430 ();
 sky130_fd_sc_hd__decap_3 PHY_1431 ();
 sky130_fd_sc_hd__decap_3 PHY_1432 ();
 sky130_fd_sc_hd__decap_3 PHY_1433 ();
 sky130_fd_sc_hd__decap_3 PHY_1434 ();
 sky130_fd_sc_hd__decap_3 PHY_1435 ();
 sky130_fd_sc_hd__decap_3 PHY_1436 ();
 sky130_fd_sc_hd__decap_3 PHY_1437 ();
 sky130_fd_sc_hd__decap_3 PHY_1438 ();
 sky130_fd_sc_hd__decap_3 PHY_1439 ();
 sky130_fd_sc_hd__decap_3 PHY_1440 ();
 sky130_fd_sc_hd__decap_3 PHY_1441 ();
 sky130_fd_sc_hd__decap_3 PHY_1442 ();
 sky130_fd_sc_hd__decap_3 PHY_1443 ();
 sky130_fd_sc_hd__decap_3 PHY_1444 ();
 sky130_fd_sc_hd__decap_3 PHY_1445 ();
 sky130_fd_sc_hd__decap_3 PHY_1446 ();
 sky130_fd_sc_hd__decap_3 PHY_1447 ();
 sky130_fd_sc_hd__decap_3 PHY_1448 ();
 sky130_fd_sc_hd__decap_3 PHY_1449 ();
 sky130_fd_sc_hd__decap_3 PHY_1450 ();
 sky130_fd_sc_hd__decap_3 PHY_1451 ();
 sky130_fd_sc_hd__decap_3 PHY_1452 ();
 sky130_fd_sc_hd__decap_3 PHY_1453 ();
 sky130_fd_sc_hd__decap_3 PHY_1454 ();
 sky130_fd_sc_hd__decap_3 PHY_1455 ();
 sky130_fd_sc_hd__decap_3 PHY_1456 ();
 sky130_fd_sc_hd__decap_3 PHY_1457 ();
 sky130_fd_sc_hd__decap_3 PHY_1458 ();
 sky130_fd_sc_hd__decap_3 PHY_1459 ();
 sky130_fd_sc_hd__decap_3 PHY_1460 ();
 sky130_fd_sc_hd__decap_3 PHY_1461 ();
 sky130_fd_sc_hd__decap_3 PHY_1462 ();
 sky130_fd_sc_hd__decap_3 PHY_1463 ();
 sky130_fd_sc_hd__decap_3 PHY_1464 ();
 sky130_fd_sc_hd__decap_3 PHY_1465 ();
 sky130_fd_sc_hd__decap_3 PHY_1466 ();
 sky130_fd_sc_hd__decap_3 PHY_1467 ();
 sky130_fd_sc_hd__decap_3 PHY_1468 ();
 sky130_fd_sc_hd__decap_3 PHY_1469 ();
 sky130_fd_sc_hd__decap_3 PHY_1470 ();
 sky130_fd_sc_hd__decap_3 PHY_1471 ();
 sky130_fd_sc_hd__decap_3 PHY_1472 ();
 sky130_fd_sc_hd__decap_3 PHY_1473 ();
 sky130_fd_sc_hd__decap_3 PHY_1474 ();
 sky130_fd_sc_hd__decap_3 PHY_1475 ();
 sky130_fd_sc_hd__decap_3 PHY_1476 ();
 sky130_fd_sc_hd__decap_3 PHY_1477 ();
 sky130_fd_sc_hd__decap_3 PHY_1478 ();
 sky130_fd_sc_hd__decap_3 PHY_1479 ();
 sky130_fd_sc_hd__decap_3 PHY_1480 ();
 sky130_fd_sc_hd__decap_3 PHY_1481 ();
 sky130_fd_sc_hd__decap_3 PHY_1482 ();
 sky130_fd_sc_hd__decap_3 PHY_1483 ();
 sky130_fd_sc_hd__decap_3 PHY_1484 ();
 sky130_fd_sc_hd__decap_3 PHY_1485 ();
 sky130_fd_sc_hd__decap_3 PHY_1486 ();
 sky130_fd_sc_hd__decap_3 PHY_1487 ();
 sky130_fd_sc_hd__decap_3 PHY_1488 ();
 sky130_fd_sc_hd__decap_3 PHY_1489 ();
 sky130_fd_sc_hd__decap_3 PHY_1490 ();
 sky130_fd_sc_hd__decap_3 PHY_1491 ();
 sky130_fd_sc_hd__decap_3 PHY_1492 ();
 sky130_fd_sc_hd__decap_3 PHY_1493 ();
 sky130_fd_sc_hd__decap_3 PHY_1494 ();
 sky130_fd_sc_hd__decap_3 PHY_1495 ();
 sky130_fd_sc_hd__decap_3 PHY_1496 ();
 sky130_fd_sc_hd__decap_3 PHY_1497 ();
 sky130_fd_sc_hd__decap_3 PHY_1498 ();
 sky130_fd_sc_hd__decap_3 PHY_1499 ();
 sky130_fd_sc_hd__decap_3 PHY_1500 ();
 sky130_fd_sc_hd__decap_3 PHY_1501 ();
 sky130_fd_sc_hd__decap_3 PHY_1502 ();
 sky130_fd_sc_hd__decap_3 PHY_1503 ();
 sky130_fd_sc_hd__decap_3 PHY_1504 ();
 sky130_fd_sc_hd__decap_3 PHY_1505 ();
 sky130_fd_sc_hd__decap_3 PHY_1506 ();
 sky130_fd_sc_hd__decap_3 PHY_1507 ();
 sky130_fd_sc_hd__decap_3 PHY_1508 ();
 sky130_fd_sc_hd__decap_3 PHY_1509 ();
 sky130_fd_sc_hd__decap_3 PHY_1510 ();
 sky130_fd_sc_hd__decap_3 PHY_1511 ();
 sky130_fd_sc_hd__decap_3 PHY_1512 ();
 sky130_fd_sc_hd__decap_3 PHY_1513 ();
 sky130_fd_sc_hd__decap_3 PHY_1514 ();
 sky130_fd_sc_hd__decap_3 PHY_1515 ();
 sky130_fd_sc_hd__decap_3 PHY_1516 ();
 sky130_fd_sc_hd__decap_3 PHY_1517 ();
 sky130_fd_sc_hd__decap_3 PHY_1518 ();
 sky130_fd_sc_hd__decap_3 PHY_1519 ();
 sky130_fd_sc_hd__decap_3 PHY_1520 ();
 sky130_fd_sc_hd__decap_3 PHY_1521 ();
 sky130_fd_sc_hd__decap_3 PHY_1522 ();
 sky130_fd_sc_hd__decap_3 PHY_1523 ();
 sky130_fd_sc_hd__decap_3 PHY_1524 ();
 sky130_fd_sc_hd__decap_3 PHY_1525 ();
 sky130_fd_sc_hd__decap_3 PHY_1526 ();
 sky130_fd_sc_hd__decap_3 PHY_1527 ();
 sky130_fd_sc_hd__decap_3 PHY_1528 ();
 sky130_fd_sc_hd__decap_3 PHY_1529 ();
 sky130_fd_sc_hd__decap_3 PHY_1530 ();
 sky130_fd_sc_hd__decap_3 PHY_1531 ();
 sky130_fd_sc_hd__decap_3 PHY_1532 ();
 sky130_fd_sc_hd__decap_3 PHY_1533 ();
 sky130_fd_sc_hd__decap_3 PHY_1534 ();
 sky130_fd_sc_hd__decap_3 PHY_1535 ();
 sky130_fd_sc_hd__decap_3 PHY_1536 ();
 sky130_fd_sc_hd__decap_3 PHY_1537 ();
 sky130_fd_sc_hd__decap_3 PHY_1538 ();
 sky130_fd_sc_hd__decap_3 PHY_1539 ();
 sky130_fd_sc_hd__decap_3 PHY_1540 ();
 sky130_fd_sc_hd__decap_3 PHY_1541 ();
 sky130_fd_sc_hd__decap_3 PHY_1542 ();
 sky130_fd_sc_hd__decap_3 PHY_1543 ();
 sky130_fd_sc_hd__decap_3 PHY_1544 ();
 sky130_fd_sc_hd__decap_3 PHY_1545 ();
 sky130_fd_sc_hd__decap_3 PHY_1546 ();
 sky130_fd_sc_hd__decap_3 PHY_1547 ();
 sky130_fd_sc_hd__decap_3 PHY_1548 ();
 sky130_fd_sc_hd__decap_3 PHY_1549 ();
 sky130_fd_sc_hd__decap_3 PHY_1550 ();
 sky130_fd_sc_hd__decap_3 PHY_1551 ();
 sky130_fd_sc_hd__decap_3 PHY_1552 ();
 sky130_fd_sc_hd__decap_3 PHY_1553 ();
 sky130_fd_sc_hd__decap_3 PHY_1554 ();
 sky130_fd_sc_hd__decap_3 PHY_1555 ();
 sky130_fd_sc_hd__decap_3 PHY_1556 ();
 sky130_fd_sc_hd__decap_3 PHY_1557 ();
 sky130_fd_sc_hd__decap_3 PHY_1558 ();
 sky130_fd_sc_hd__decap_3 PHY_1559 ();
 sky130_fd_sc_hd__decap_3 PHY_1560 ();
 sky130_fd_sc_hd__decap_3 PHY_1561 ();
 sky130_fd_sc_hd__decap_3 PHY_1562 ();
 sky130_fd_sc_hd__decap_3 PHY_1563 ();
 sky130_fd_sc_hd__decap_3 PHY_1564 ();
 sky130_fd_sc_hd__decap_3 PHY_1565 ();
 sky130_fd_sc_hd__decap_3 PHY_1566 ();
 sky130_fd_sc_hd__decap_3 PHY_1567 ();
 sky130_fd_sc_hd__decap_3 PHY_1568 ();
 sky130_fd_sc_hd__decap_3 PHY_1569 ();
 sky130_fd_sc_hd__decap_3 PHY_1570 ();
 sky130_fd_sc_hd__decap_3 PHY_1571 ();
 sky130_fd_sc_hd__decap_3 PHY_1572 ();
 sky130_fd_sc_hd__decap_3 PHY_1573 ();
 sky130_fd_sc_hd__decap_3 PHY_1574 ();
 sky130_fd_sc_hd__decap_3 PHY_1575 ();
 sky130_fd_sc_hd__decap_3 PHY_1576 ();
 sky130_fd_sc_hd__decap_3 PHY_1577 ();
 sky130_fd_sc_hd__decap_3 PHY_1578 ();
 sky130_fd_sc_hd__decap_3 PHY_1579 ();
 sky130_fd_sc_hd__decap_3 PHY_1580 ();
 sky130_fd_sc_hd__decap_3 PHY_1581 ();
 sky130_fd_sc_hd__decap_3 PHY_1582 ();
 sky130_fd_sc_hd__decap_3 PHY_1583 ();
 sky130_fd_sc_hd__decap_3 PHY_1584 ();
 sky130_fd_sc_hd__decap_3 PHY_1585 ();
 sky130_fd_sc_hd__decap_3 PHY_1586 ();
 sky130_fd_sc_hd__decap_3 PHY_1587 ();
 sky130_fd_sc_hd__decap_3 PHY_1588 ();
 sky130_fd_sc_hd__decap_3 PHY_1589 ();
 sky130_fd_sc_hd__decap_3 PHY_1590 ();
 sky130_fd_sc_hd__decap_3 PHY_1591 ();
 sky130_fd_sc_hd__decap_3 PHY_1592 ();
 sky130_fd_sc_hd__decap_3 PHY_1593 ();
 sky130_fd_sc_hd__decap_3 PHY_1594 ();
 sky130_fd_sc_hd__decap_3 PHY_1595 ();
 sky130_fd_sc_hd__decap_3 PHY_1596 ();
 sky130_fd_sc_hd__decap_3 PHY_1597 ();
 sky130_fd_sc_hd__decap_3 PHY_1598 ();
 sky130_fd_sc_hd__decap_3 PHY_1599 ();
 sky130_fd_sc_hd__decap_3 PHY_1600 ();
 sky130_fd_sc_hd__decap_3 PHY_1601 ();
 sky130_fd_sc_hd__decap_3 PHY_1602 ();
 sky130_fd_sc_hd__decap_3 PHY_1603 ();
 sky130_fd_sc_hd__decap_3 PHY_1604 ();
 sky130_fd_sc_hd__decap_3 PHY_1605 ();
 sky130_fd_sc_hd__decap_3 PHY_1606 ();
 sky130_fd_sc_hd__decap_3 PHY_1607 ();
 sky130_fd_sc_hd__decap_3 PHY_1608 ();
 sky130_fd_sc_hd__decap_3 PHY_1609 ();
 sky130_fd_sc_hd__decap_3 PHY_1610 ();
 sky130_fd_sc_hd__decap_3 PHY_1611 ();
 sky130_fd_sc_hd__decap_3 PHY_1612 ();
 sky130_fd_sc_hd__decap_3 PHY_1613 ();
 sky130_fd_sc_hd__decap_3 PHY_1614 ();
 sky130_fd_sc_hd__decap_3 PHY_1615 ();
 sky130_fd_sc_hd__decap_3 PHY_1616 ();
 sky130_fd_sc_hd__decap_3 PHY_1617 ();
 sky130_fd_sc_hd__decap_3 PHY_1618 ();
 sky130_fd_sc_hd__decap_3 PHY_1619 ();
 sky130_fd_sc_hd__decap_3 PHY_1620 ();
 sky130_fd_sc_hd__decap_3 PHY_1621 ();
 sky130_fd_sc_hd__decap_3 PHY_1622 ();
 sky130_fd_sc_hd__decap_3 PHY_1623 ();
 sky130_fd_sc_hd__decap_3 PHY_1624 ();
 sky130_fd_sc_hd__decap_3 PHY_1625 ();
 sky130_fd_sc_hd__decap_3 PHY_1626 ();
 sky130_fd_sc_hd__decap_3 PHY_1627 ();
 sky130_fd_sc_hd__decap_3 PHY_1628 ();
 sky130_fd_sc_hd__decap_3 PHY_1629 ();
 sky130_fd_sc_hd__decap_3 PHY_1630 ();
 sky130_fd_sc_hd__decap_3 PHY_1631 ();
 sky130_fd_sc_hd__decap_3 PHY_1632 ();
 sky130_fd_sc_hd__decap_3 PHY_1633 ();
 sky130_fd_sc_hd__decap_3 PHY_1634 ();
 sky130_fd_sc_hd__decap_3 PHY_1635 ();
 sky130_fd_sc_hd__decap_3 PHY_1636 ();
 sky130_fd_sc_hd__decap_3 PHY_1637 ();
 sky130_fd_sc_hd__decap_3 PHY_1638 ();
 sky130_fd_sc_hd__decap_3 PHY_1639 ();
 sky130_fd_sc_hd__decap_3 PHY_1640 ();
 sky130_fd_sc_hd__decap_3 PHY_1641 ();
 sky130_fd_sc_hd__decap_3 PHY_1642 ();
 sky130_fd_sc_hd__decap_3 PHY_1643 ();
 sky130_fd_sc_hd__decap_3 PHY_1644 ();
 sky130_fd_sc_hd__decap_3 PHY_1645 ();
 sky130_fd_sc_hd__decap_3 PHY_1646 ();
 sky130_fd_sc_hd__decap_3 PHY_1647 ();
 sky130_fd_sc_hd__decap_3 PHY_1648 ();
 sky130_fd_sc_hd__decap_3 PHY_1649 ();
 sky130_fd_sc_hd__decap_3 PHY_1650 ();
 sky130_fd_sc_hd__decap_3 PHY_1651 ();
 sky130_fd_sc_hd__decap_3 PHY_1652 ();
 sky130_fd_sc_hd__decap_3 PHY_1653 ();
 sky130_fd_sc_hd__decap_3 PHY_1654 ();
 sky130_fd_sc_hd__decap_3 PHY_1655 ();
 sky130_fd_sc_hd__decap_3 PHY_1656 ();
 sky130_fd_sc_hd__decap_3 PHY_1657 ();
 sky130_fd_sc_hd__decap_3 PHY_1658 ();
 sky130_fd_sc_hd__decap_3 PHY_1659 ();
 sky130_fd_sc_hd__decap_3 PHY_1660 ();
 sky130_fd_sc_hd__decap_3 PHY_1661 ();
 sky130_fd_sc_hd__decap_3 PHY_1662 ();
 sky130_fd_sc_hd__decap_3 PHY_1663 ();
 sky130_fd_sc_hd__decap_3 PHY_1664 ();
 sky130_fd_sc_hd__decap_3 PHY_1665 ();
 sky130_fd_sc_hd__decap_3 PHY_1666 ();
 sky130_fd_sc_hd__decap_3 PHY_1667 ();
 sky130_fd_sc_hd__decap_3 PHY_1668 ();
 sky130_fd_sc_hd__decap_3 PHY_1669 ();
 sky130_fd_sc_hd__decap_3 PHY_1670 ();
 sky130_fd_sc_hd__decap_3 PHY_1671 ();
 sky130_fd_sc_hd__decap_3 PHY_1672 ();
 sky130_fd_sc_hd__decap_3 PHY_1673 ();
 sky130_fd_sc_hd__decap_3 PHY_1674 ();
 sky130_fd_sc_hd__decap_3 PHY_1675 ();
 sky130_fd_sc_hd__decap_3 PHY_1676 ();
 sky130_fd_sc_hd__decap_3 PHY_1677 ();
 sky130_fd_sc_hd__decap_3 PHY_1678 ();
 sky130_fd_sc_hd__decap_3 PHY_1679 ();
 sky130_fd_sc_hd__decap_3 PHY_1680 ();
 sky130_fd_sc_hd__decap_3 PHY_1681 ();
 sky130_fd_sc_hd__decap_3 PHY_1682 ();
 sky130_fd_sc_hd__decap_3 PHY_1683 ();
 sky130_fd_sc_hd__decap_3 PHY_1684 ();
 sky130_fd_sc_hd__decap_3 PHY_1685 ();
 sky130_fd_sc_hd__decap_3 PHY_1686 ();
 sky130_fd_sc_hd__decap_3 PHY_1687 ();
 sky130_fd_sc_hd__decap_3 PHY_1688 ();
 sky130_fd_sc_hd__decap_3 PHY_1689 ();
 sky130_fd_sc_hd__decap_3 PHY_1690 ();
 sky130_fd_sc_hd__decap_3 PHY_1691 ();
 sky130_fd_sc_hd__decap_3 PHY_1692 ();
 sky130_fd_sc_hd__decap_3 PHY_1693 ();
 sky130_fd_sc_hd__decap_3 PHY_1694 ();
 sky130_fd_sc_hd__decap_3 PHY_1695 ();
 sky130_fd_sc_hd__decap_3 PHY_1696 ();
 sky130_fd_sc_hd__decap_3 PHY_1697 ();
 sky130_fd_sc_hd__decap_3 PHY_1698 ();
 sky130_fd_sc_hd__decap_3 PHY_1699 ();
 sky130_fd_sc_hd__decap_3 PHY_1700 ();
 sky130_fd_sc_hd__decap_3 PHY_1701 ();
 sky130_fd_sc_hd__decap_3 PHY_1702 ();
 sky130_fd_sc_hd__decap_3 PHY_1703 ();
 sky130_fd_sc_hd__decap_3 PHY_1704 ();
 sky130_fd_sc_hd__decap_3 PHY_1705 ();
 sky130_fd_sc_hd__decap_3 PHY_1706 ();
 sky130_fd_sc_hd__decap_3 PHY_1707 ();
 sky130_fd_sc_hd__decap_3 PHY_1708 ();
 sky130_fd_sc_hd__decap_3 PHY_1709 ();
 sky130_fd_sc_hd__decap_3 PHY_1710 ();
 sky130_fd_sc_hd__decap_3 PHY_1711 ();
 sky130_fd_sc_hd__decap_3 PHY_1712 ();
 sky130_fd_sc_hd__decap_3 PHY_1713 ();
 sky130_fd_sc_hd__decap_3 PHY_1714 ();
 sky130_fd_sc_hd__decap_3 PHY_1715 ();
 sky130_fd_sc_hd__decap_3 PHY_1716 ();
 sky130_fd_sc_hd__decap_3 PHY_1717 ();
 sky130_fd_sc_hd__decap_3 PHY_1718 ();
 sky130_fd_sc_hd__decap_3 PHY_1719 ();
 sky130_fd_sc_hd__decap_3 PHY_1720 ();
 sky130_fd_sc_hd__decap_3 PHY_1721 ();
 sky130_fd_sc_hd__decap_3 PHY_1722 ();
 sky130_fd_sc_hd__decap_3 PHY_1723 ();
 sky130_fd_sc_hd__decap_3 PHY_1724 ();
 sky130_fd_sc_hd__decap_3 PHY_1725 ();
 sky130_fd_sc_hd__decap_3 PHY_1726 ();
 sky130_fd_sc_hd__decap_3 PHY_1727 ();
 sky130_fd_sc_hd__decap_3 PHY_1728 ();
 sky130_fd_sc_hd__decap_3 PHY_1729 ();
 sky130_fd_sc_hd__decap_3 PHY_1730 ();
 sky130_fd_sc_hd__decap_3 PHY_1731 ();
 sky130_fd_sc_hd__decap_3 PHY_1732 ();
 sky130_fd_sc_hd__decap_3 PHY_1733 ();
 sky130_fd_sc_hd__decap_3 PHY_1734 ();
 sky130_fd_sc_hd__decap_3 PHY_1735 ();
 sky130_fd_sc_hd__decap_3 PHY_1736 ();
 sky130_fd_sc_hd__decap_3 PHY_1737 ();
 sky130_fd_sc_hd__decap_3 PHY_1738 ();
 sky130_fd_sc_hd__decap_3 PHY_1739 ();
 sky130_fd_sc_hd__decap_3 PHY_1740 ();
 sky130_fd_sc_hd__decap_3 PHY_1741 ();
 sky130_fd_sc_hd__decap_3 PHY_1742 ();
 sky130_fd_sc_hd__decap_3 PHY_1743 ();
 sky130_fd_sc_hd__decap_3 PHY_1744 ();
 sky130_fd_sc_hd__decap_3 PHY_1745 ();
 sky130_fd_sc_hd__decap_3 PHY_1746 ();
 sky130_fd_sc_hd__decap_3 PHY_1747 ();
 sky130_fd_sc_hd__decap_3 PHY_1748 ();
 sky130_fd_sc_hd__decap_3 PHY_1749 ();
 sky130_fd_sc_hd__decap_3 PHY_1750 ();
 sky130_fd_sc_hd__decap_3 PHY_1751 ();
 sky130_fd_sc_hd__decap_3 PHY_1752 ();
 sky130_fd_sc_hd__decap_3 PHY_1753 ();
 sky130_fd_sc_hd__decap_3 PHY_1754 ();
 sky130_fd_sc_hd__decap_3 PHY_1755 ();
 sky130_fd_sc_hd__decap_3 PHY_1756 ();
 sky130_fd_sc_hd__decap_3 PHY_1757 ();
 sky130_fd_sc_hd__decap_3 PHY_1758 ();
 sky130_fd_sc_hd__decap_3 PHY_1759 ();
 sky130_fd_sc_hd__decap_3 PHY_1760 ();
 sky130_fd_sc_hd__decap_3 PHY_1761 ();
 sky130_fd_sc_hd__decap_3 PHY_1762 ();
 sky130_fd_sc_hd__decap_3 PHY_1763 ();
 sky130_fd_sc_hd__decap_3 PHY_1764 ();
 sky130_fd_sc_hd__decap_3 PHY_1765 ();
 sky130_fd_sc_hd__decap_3 PHY_1766 ();
 sky130_fd_sc_hd__decap_3 PHY_1767 ();
 sky130_fd_sc_hd__decap_3 PHY_1768 ();
 sky130_fd_sc_hd__decap_3 PHY_1769 ();
 sky130_fd_sc_hd__decap_3 PHY_1770 ();
 sky130_fd_sc_hd__decap_3 PHY_1771 ();
 sky130_fd_sc_hd__decap_3 PHY_1772 ();
 sky130_fd_sc_hd__decap_3 PHY_1773 ();
 sky130_fd_sc_hd__decap_3 PHY_1774 ();
 sky130_fd_sc_hd__decap_3 PHY_1775 ();
 sky130_fd_sc_hd__decap_3 PHY_1776 ();
 sky130_fd_sc_hd__decap_3 PHY_1777 ();
 sky130_fd_sc_hd__decap_3 PHY_1778 ();
 sky130_fd_sc_hd__decap_3 PHY_1779 ();
 sky130_fd_sc_hd__decap_3 PHY_1780 ();
 sky130_fd_sc_hd__decap_3 PHY_1781 ();
 sky130_fd_sc_hd__decap_3 PHY_1782 ();
 sky130_fd_sc_hd__decap_3 PHY_1783 ();
 sky130_fd_sc_hd__decap_3 PHY_1784 ();
 sky130_fd_sc_hd__decap_3 PHY_1785 ();
 sky130_fd_sc_hd__decap_3 PHY_1786 ();
 sky130_fd_sc_hd__decap_3 PHY_1787 ();
 sky130_fd_sc_hd__decap_3 PHY_1788 ();
 sky130_fd_sc_hd__decap_3 PHY_1789 ();
 sky130_fd_sc_hd__decap_3 PHY_1790 ();
 sky130_fd_sc_hd__decap_3 PHY_1791 ();
 sky130_fd_sc_hd__decap_3 PHY_1792 ();
 sky130_fd_sc_hd__decap_3 PHY_1793 ();
 sky130_fd_sc_hd__decap_3 PHY_1794 ();
 sky130_fd_sc_hd__decap_3 PHY_1795 ();
 sky130_fd_sc_hd__decap_3 PHY_1796 ();
 sky130_fd_sc_hd__decap_3 PHY_1797 ();
 sky130_fd_sc_hd__decap_3 PHY_1798 ();
 sky130_fd_sc_hd__decap_3 PHY_1799 ();
 sky130_fd_sc_hd__decap_3 PHY_1800 ();
 sky130_fd_sc_hd__decap_3 PHY_1801 ();
 sky130_fd_sc_hd__decap_3 PHY_1802 ();
 sky130_fd_sc_hd__decap_3 PHY_1803 ();
 sky130_fd_sc_hd__decap_3 PHY_1804 ();
 sky130_fd_sc_hd__decap_3 PHY_1805 ();
 sky130_fd_sc_hd__decap_3 PHY_1806 ();
 sky130_fd_sc_hd__decap_3 PHY_1807 ();
 sky130_fd_sc_hd__decap_3 PHY_1808 ();
 sky130_fd_sc_hd__decap_3 PHY_1809 ();
 sky130_fd_sc_hd__decap_3 PHY_1810 ();
 sky130_fd_sc_hd__decap_3 PHY_1811 ();
 sky130_fd_sc_hd__decap_3 PHY_1812 ();
 sky130_fd_sc_hd__decap_3 PHY_1813 ();
 sky130_fd_sc_hd__decap_3 PHY_1814 ();
 sky130_fd_sc_hd__decap_3 PHY_1815 ();
 sky130_fd_sc_hd__decap_3 PHY_1816 ();
 sky130_fd_sc_hd__decap_3 PHY_1817 ();
 sky130_fd_sc_hd__decap_3 PHY_1818 ();
 sky130_fd_sc_hd__decap_3 PHY_1819 ();
 sky130_fd_sc_hd__decap_3 PHY_1820 ();
 sky130_fd_sc_hd__decap_3 PHY_1821 ();
 sky130_fd_sc_hd__decap_3 PHY_1822 ();
 sky130_fd_sc_hd__decap_3 PHY_1823 ();
 sky130_fd_sc_hd__decap_3 PHY_1824 ();
 sky130_fd_sc_hd__decap_3 PHY_1825 ();
 sky130_fd_sc_hd__decap_3 PHY_1826 ();
 sky130_fd_sc_hd__decap_3 PHY_1827 ();
 sky130_fd_sc_hd__decap_3 PHY_1828 ();
 sky130_fd_sc_hd__decap_3 PHY_1829 ();
 sky130_fd_sc_hd__decap_3 PHY_1830 ();
 sky130_fd_sc_hd__decap_3 PHY_1831 ();
 sky130_fd_sc_hd__decap_3 PHY_1832 ();
 sky130_fd_sc_hd__decap_3 PHY_1833 ();
 sky130_fd_sc_hd__decap_3 PHY_1834 ();
 sky130_fd_sc_hd__decap_3 PHY_1835 ();
 sky130_fd_sc_hd__decap_3 PHY_1836 ();
 sky130_fd_sc_hd__decap_3 PHY_1837 ();
 sky130_fd_sc_hd__decap_3 PHY_1838 ();
 sky130_fd_sc_hd__decap_3 PHY_1839 ();
 sky130_fd_sc_hd__decap_3 PHY_1840 ();
 sky130_fd_sc_hd__decap_3 PHY_1841 ();
 sky130_fd_sc_hd__decap_3 PHY_1842 ();
 sky130_fd_sc_hd__decap_3 PHY_1843 ();
 sky130_fd_sc_hd__decap_3 PHY_1844 ();
 sky130_fd_sc_hd__decap_3 PHY_1845 ();
 sky130_fd_sc_hd__decap_3 PHY_1846 ();
 sky130_fd_sc_hd__decap_3 PHY_1847 ();
 sky130_fd_sc_hd__decap_3 PHY_1848 ();
 sky130_fd_sc_hd__decap_3 PHY_1849 ();
 sky130_fd_sc_hd__decap_3 PHY_1850 ();
 sky130_fd_sc_hd__decap_3 PHY_1851 ();
 sky130_fd_sc_hd__decap_3 PHY_1852 ();
 sky130_fd_sc_hd__decap_3 PHY_1853 ();
 sky130_fd_sc_hd__decap_3 PHY_1854 ();
 sky130_fd_sc_hd__decap_3 PHY_1855 ();
 sky130_fd_sc_hd__decap_3 PHY_1856 ();
 sky130_fd_sc_hd__decap_3 PHY_1857 ();
 sky130_fd_sc_hd__decap_3 PHY_1858 ();
 sky130_fd_sc_hd__decap_3 PHY_1859 ();
 sky130_fd_sc_hd__decap_3 PHY_1860 ();
 sky130_fd_sc_hd__decap_3 PHY_1861 ();
 sky130_fd_sc_hd__decap_3 PHY_1862 ();
 sky130_fd_sc_hd__decap_3 PHY_1863 ();
 sky130_fd_sc_hd__decap_3 PHY_1864 ();
 sky130_fd_sc_hd__decap_3 PHY_1865 ();
 sky130_fd_sc_hd__decap_3 PHY_1866 ();
 sky130_fd_sc_hd__decap_3 PHY_1867 ();
 sky130_fd_sc_hd__decap_3 PHY_1868 ();
 sky130_fd_sc_hd__decap_3 PHY_1869 ();
 sky130_fd_sc_hd__decap_3 PHY_1870 ();
 sky130_fd_sc_hd__decap_3 PHY_1871 ();
 sky130_fd_sc_hd__decap_3 PHY_1872 ();
 sky130_fd_sc_hd__decap_3 PHY_1873 ();
 sky130_fd_sc_hd__decap_3 PHY_1874 ();
 sky130_fd_sc_hd__decap_3 PHY_1875 ();
 sky130_fd_sc_hd__decap_3 PHY_1876 ();
 sky130_fd_sc_hd__decap_3 PHY_1877 ();
 sky130_fd_sc_hd__decap_3 PHY_1878 ();
 sky130_fd_sc_hd__decap_3 PHY_1879 ();
 sky130_fd_sc_hd__decap_3 PHY_1880 ();
 sky130_fd_sc_hd__decap_3 PHY_1881 ();
 sky130_fd_sc_hd__decap_3 PHY_1882 ();
 sky130_fd_sc_hd__decap_3 PHY_1883 ();
 sky130_fd_sc_hd__decap_3 PHY_1884 ();
 sky130_fd_sc_hd__decap_3 PHY_1885 ();
 sky130_fd_sc_hd__decap_3 PHY_1886 ();
 sky130_fd_sc_hd__decap_3 PHY_1887 ();
 sky130_fd_sc_hd__decap_3 PHY_1888 ();
 sky130_fd_sc_hd__decap_3 PHY_1889 ();
 sky130_fd_sc_hd__decap_3 PHY_1890 ();
 sky130_fd_sc_hd__decap_3 PHY_1891 ();
 sky130_fd_sc_hd__decap_3 PHY_1892 ();
 sky130_fd_sc_hd__decap_3 PHY_1893 ();
 sky130_fd_sc_hd__decap_3 PHY_1894 ();
 sky130_fd_sc_hd__decap_3 PHY_1895 ();
 sky130_fd_sc_hd__decap_3 PHY_1896 ();
 sky130_fd_sc_hd__decap_3 PHY_1897 ();
 sky130_fd_sc_hd__decap_3 PHY_1898 ();
 sky130_fd_sc_hd__decap_3 PHY_1899 ();
 sky130_fd_sc_hd__decap_3 PHY_1900 ();
 sky130_fd_sc_hd__decap_3 PHY_1901 ();
 sky130_fd_sc_hd__decap_3 PHY_1902 ();
 sky130_fd_sc_hd__decap_3 PHY_1903 ();
 sky130_fd_sc_hd__decap_3 PHY_1904 ();
 sky130_fd_sc_hd__decap_3 PHY_1905 ();
 sky130_fd_sc_hd__decap_3 PHY_1906 ();
 sky130_fd_sc_hd__decap_3 PHY_1907 ();
 sky130_fd_sc_hd__decap_3 PHY_1908 ();
 sky130_fd_sc_hd__decap_3 PHY_1909 ();
 sky130_fd_sc_hd__decap_3 PHY_1910 ();
 sky130_fd_sc_hd__decap_3 PHY_1911 ();
 sky130_fd_sc_hd__decap_3 PHY_1912 ();
 sky130_fd_sc_hd__decap_3 PHY_1913 ();
 sky130_fd_sc_hd__decap_3 PHY_1914 ();
 sky130_fd_sc_hd__decap_3 PHY_1915 ();
 sky130_fd_sc_hd__decap_3 PHY_1916 ();
 sky130_fd_sc_hd__decap_3 PHY_1917 ();
 sky130_fd_sc_hd__decap_3 PHY_1918 ();
 sky130_fd_sc_hd__decap_3 PHY_1919 ();
 sky130_fd_sc_hd__decap_3 PHY_1920 ();
 sky130_fd_sc_hd__decap_3 PHY_1921 ();
 sky130_fd_sc_hd__decap_3 PHY_1922 ();
 sky130_fd_sc_hd__decap_3 PHY_1923 ();
 sky130_fd_sc_hd__decap_3 PHY_1924 ();
 sky130_fd_sc_hd__decap_3 PHY_1925 ();
 sky130_fd_sc_hd__decap_3 PHY_1926 ();
 sky130_fd_sc_hd__decap_3 PHY_1927 ();
 sky130_fd_sc_hd__decap_3 PHY_1928 ();
 sky130_fd_sc_hd__decap_3 PHY_1929 ();
 sky130_fd_sc_hd__decap_3 PHY_1930 ();
 sky130_fd_sc_hd__decap_3 PHY_1931 ();
 sky130_fd_sc_hd__decap_3 PHY_1932 ();
 sky130_fd_sc_hd__decap_3 PHY_1933 ();
 sky130_fd_sc_hd__decap_3 PHY_1934 ();
 sky130_fd_sc_hd__decap_3 PHY_1935 ();
 sky130_fd_sc_hd__decap_3 PHY_1936 ();
 sky130_fd_sc_hd__decap_3 PHY_1937 ();
 sky130_fd_sc_hd__decap_3 PHY_1938 ();
 sky130_fd_sc_hd__decap_3 PHY_1939 ();
 sky130_fd_sc_hd__decap_3 PHY_1940 ();
 sky130_fd_sc_hd__decap_3 PHY_1941 ();
 sky130_fd_sc_hd__decap_3 PHY_1942 ();
 sky130_fd_sc_hd__decap_3 PHY_1943 ();
 sky130_fd_sc_hd__decap_3 PHY_1944 ();
 sky130_fd_sc_hd__decap_3 PHY_1945 ();
 sky130_fd_sc_hd__decap_3 PHY_1946 ();
 sky130_fd_sc_hd__decap_3 PHY_1947 ();
 sky130_fd_sc_hd__decap_3 PHY_1948 ();
 sky130_fd_sc_hd__decap_3 PHY_1949 ();
 sky130_fd_sc_hd__decap_3 PHY_1950 ();
 sky130_fd_sc_hd__decap_3 PHY_1951 ();
 sky130_fd_sc_hd__decap_3 PHY_1952 ();
 sky130_fd_sc_hd__decap_3 PHY_1953 ();
 sky130_fd_sc_hd__decap_3 PHY_1954 ();
 sky130_fd_sc_hd__decap_3 PHY_1955 ();
 sky130_fd_sc_hd__decap_3 PHY_1956 ();
 sky130_fd_sc_hd__decap_3 PHY_1957 ();
 sky130_fd_sc_hd__decap_3 PHY_1958 ();
 sky130_fd_sc_hd__decap_3 PHY_1959 ();
 sky130_fd_sc_hd__decap_3 PHY_1960 ();
 sky130_fd_sc_hd__decap_3 PHY_1961 ();
 sky130_fd_sc_hd__decap_3 PHY_1962 ();
 sky130_fd_sc_hd__decap_3 PHY_1963 ();
 sky130_fd_sc_hd__decap_3 PHY_1964 ();
 sky130_fd_sc_hd__decap_3 PHY_1965 ();
 sky130_fd_sc_hd__decap_3 PHY_1966 ();
 sky130_fd_sc_hd__decap_3 PHY_1967 ();
 sky130_fd_sc_hd__decap_3 PHY_1968 ();
 sky130_fd_sc_hd__decap_3 PHY_1969 ();
 sky130_fd_sc_hd__decap_3 PHY_1970 ();
 sky130_fd_sc_hd__decap_3 PHY_1971 ();
 sky130_fd_sc_hd__decap_3 PHY_1972 ();
 sky130_fd_sc_hd__decap_3 PHY_1973 ();
 sky130_fd_sc_hd__decap_3 PHY_1974 ();
 sky130_fd_sc_hd__decap_3 PHY_1975 ();
 sky130_fd_sc_hd__decap_3 PHY_1976 ();
 sky130_fd_sc_hd__decap_3 PHY_1977 ();
 sky130_fd_sc_hd__decap_3 PHY_1978 ();
 sky130_fd_sc_hd__decap_3 PHY_1979 ();
 sky130_fd_sc_hd__decap_3 PHY_1980 ();
 sky130_fd_sc_hd__decap_3 PHY_1981 ();
 sky130_fd_sc_hd__decap_3 PHY_1982 ();
 sky130_fd_sc_hd__decap_3 PHY_1983 ();
 sky130_fd_sc_hd__decap_3 PHY_1984 ();
 sky130_fd_sc_hd__decap_3 PHY_1985 ();
 sky130_fd_sc_hd__decap_3 PHY_1986 ();
 sky130_fd_sc_hd__decap_3 PHY_1987 ();
 sky130_fd_sc_hd__decap_3 PHY_1988 ();
 sky130_fd_sc_hd__decap_3 PHY_1989 ();
 sky130_fd_sc_hd__decap_3 PHY_1990 ();
 sky130_fd_sc_hd__decap_3 PHY_1991 ();
 sky130_fd_sc_hd__decap_3 PHY_1992 ();
 sky130_fd_sc_hd__decap_3 PHY_1993 ();
 sky130_fd_sc_hd__decap_3 PHY_1994 ();
 sky130_fd_sc_hd__decap_3 PHY_1995 ();
 sky130_fd_sc_hd__decap_3 PHY_1996 ();
 sky130_fd_sc_hd__decap_3 PHY_1997 ();
 sky130_fd_sc_hd__decap_3 PHY_1998 ();
 sky130_fd_sc_hd__decap_3 PHY_1999 ();
 sky130_fd_sc_hd__decap_3 PHY_2000 ();
 sky130_fd_sc_hd__decap_3 PHY_2001 ();
 sky130_fd_sc_hd__decap_3 PHY_2002 ();
 sky130_fd_sc_hd__decap_3 PHY_2003 ();
 sky130_fd_sc_hd__decap_3 PHY_2004 ();
 sky130_fd_sc_hd__decap_3 PHY_2005 ();
 sky130_fd_sc_hd__decap_3 PHY_2006 ();
 sky130_fd_sc_hd__decap_3 PHY_2007 ();
 sky130_fd_sc_hd__decap_3 PHY_2008 ();
 sky130_fd_sc_hd__decap_3 PHY_2009 ();
 sky130_fd_sc_hd__decap_3 PHY_2010 ();
 sky130_fd_sc_hd__decap_3 PHY_2011 ();
 sky130_fd_sc_hd__decap_3 PHY_2012 ();
 sky130_fd_sc_hd__decap_3 PHY_2013 ();
 sky130_fd_sc_hd__decap_3 PHY_2014 ();
 sky130_fd_sc_hd__decap_3 PHY_2015 ();
 sky130_fd_sc_hd__decap_3 PHY_2016 ();
 sky130_fd_sc_hd__decap_3 PHY_2017 ();
 sky130_fd_sc_hd__decap_3 PHY_2018 ();
 sky130_fd_sc_hd__decap_3 PHY_2019 ();
 sky130_fd_sc_hd__decap_3 PHY_2020 ();
 sky130_fd_sc_hd__decap_3 PHY_2021 ();
 sky130_fd_sc_hd__decap_3 PHY_2022 ();
 sky130_fd_sc_hd__decap_3 PHY_2023 ();
 sky130_fd_sc_hd__decap_3 PHY_2024 ();
 sky130_fd_sc_hd__decap_3 PHY_2025 ();
 sky130_fd_sc_hd__decap_3 PHY_2026 ();
 sky130_fd_sc_hd__decap_3 PHY_2027 ();
 sky130_fd_sc_hd__decap_3 PHY_2028 ();
 sky130_fd_sc_hd__decap_3 PHY_2029 ();
 sky130_fd_sc_hd__decap_3 PHY_2030 ();
 sky130_fd_sc_hd__decap_3 PHY_2031 ();
 sky130_fd_sc_hd__decap_3 PHY_2032 ();
 sky130_fd_sc_hd__decap_3 PHY_2033 ();
 sky130_fd_sc_hd__decap_3 PHY_2034 ();
 sky130_fd_sc_hd__decap_3 PHY_2035 ();
 sky130_fd_sc_hd__decap_3 PHY_2036 ();
 sky130_fd_sc_hd__decap_3 PHY_2037 ();
 sky130_fd_sc_hd__decap_3 PHY_2038 ();
 sky130_fd_sc_hd__decap_3 PHY_2039 ();
 sky130_fd_sc_hd__decap_3 PHY_2040 ();
 sky130_fd_sc_hd__decap_3 PHY_2041 ();
 sky130_fd_sc_hd__decap_3 PHY_2042 ();
 sky130_fd_sc_hd__decap_3 PHY_2043 ();
 sky130_fd_sc_hd__decap_3 PHY_2044 ();
 sky130_fd_sc_hd__decap_3 PHY_2045 ();
 sky130_fd_sc_hd__decap_3 PHY_2046 ();
 sky130_fd_sc_hd__decap_3 PHY_2047 ();
 sky130_fd_sc_hd__decap_3 PHY_2048 ();
 sky130_fd_sc_hd__decap_3 PHY_2049 ();
 sky130_fd_sc_hd__decap_3 PHY_2050 ();
 sky130_fd_sc_hd__decap_3 PHY_2051 ();
 sky130_fd_sc_hd__decap_3 PHY_2052 ();
 sky130_fd_sc_hd__decap_3 PHY_2053 ();
 sky130_fd_sc_hd__decap_3 PHY_2054 ();
 sky130_fd_sc_hd__decap_3 PHY_2055 ();
 sky130_fd_sc_hd__decap_3 PHY_2056 ();
 sky130_fd_sc_hd__decap_3 PHY_2057 ();
 sky130_fd_sc_hd__decap_3 PHY_2058 ();
 sky130_fd_sc_hd__decap_3 PHY_2059 ();
 sky130_fd_sc_hd__decap_3 PHY_2060 ();
 sky130_fd_sc_hd__decap_3 PHY_2061 ();
 sky130_fd_sc_hd__decap_3 PHY_2062 ();
 sky130_fd_sc_hd__decap_3 PHY_2063 ();
 sky130_fd_sc_hd__decap_3 PHY_2064 ();
 sky130_fd_sc_hd__decap_3 PHY_2065 ();
 sky130_fd_sc_hd__decap_3 PHY_2066 ();
 sky130_fd_sc_hd__decap_3 PHY_2067 ();
 sky130_fd_sc_hd__decap_3 PHY_2068 ();
 sky130_fd_sc_hd__decap_3 PHY_2069 ();
 sky130_fd_sc_hd__decap_3 PHY_2070 ();
 sky130_fd_sc_hd__decap_3 PHY_2071 ();
 sky130_fd_sc_hd__decap_3 PHY_2072 ();
 sky130_fd_sc_hd__decap_3 PHY_2073 ();
 sky130_fd_sc_hd__decap_3 PHY_2074 ();
 sky130_fd_sc_hd__decap_3 PHY_2075 ();
 sky130_fd_sc_hd__decap_3 PHY_2076 ();
 sky130_fd_sc_hd__decap_3 PHY_2077 ();
 sky130_fd_sc_hd__decap_3 PHY_2078 ();
 sky130_fd_sc_hd__decap_3 PHY_2079 ();
 sky130_fd_sc_hd__decap_3 PHY_2080 ();
 sky130_fd_sc_hd__decap_3 PHY_2081 ();
 sky130_fd_sc_hd__decap_3 PHY_2082 ();
 sky130_fd_sc_hd__decap_3 PHY_2083 ();
 sky130_fd_sc_hd__decap_3 PHY_2084 ();
 sky130_fd_sc_hd__decap_3 PHY_2085 ();
 sky130_fd_sc_hd__decap_3 PHY_2086 ();
 sky130_fd_sc_hd__decap_3 PHY_2087 ();
 sky130_fd_sc_hd__decap_3 PHY_2088 ();
 sky130_fd_sc_hd__decap_3 PHY_2089 ();
 sky130_fd_sc_hd__decap_3 PHY_2090 ();
 sky130_fd_sc_hd__decap_3 PHY_2091 ();
 sky130_fd_sc_hd__decap_3 PHY_2092 ();
 sky130_fd_sc_hd__decap_3 PHY_2093 ();
 sky130_fd_sc_hd__decap_3 PHY_2094 ();
 sky130_fd_sc_hd__decap_3 PHY_2095 ();
 sky130_fd_sc_hd__decap_3 PHY_2096 ();
 sky130_fd_sc_hd__decap_3 PHY_2097 ();
 sky130_fd_sc_hd__decap_3 PHY_2098 ();
 sky130_fd_sc_hd__decap_3 PHY_2099 ();
 sky130_fd_sc_hd__decap_3 PHY_2100 ();
 sky130_fd_sc_hd__decap_3 PHY_2101 ();
 sky130_fd_sc_hd__decap_3 PHY_2102 ();
 sky130_fd_sc_hd__decap_3 PHY_2103 ();
 sky130_fd_sc_hd__decap_3 PHY_2104 ();
 sky130_fd_sc_hd__decap_3 PHY_2105 ();
 sky130_fd_sc_hd__decap_3 PHY_2106 ();
 sky130_fd_sc_hd__decap_3 PHY_2107 ();
 sky130_fd_sc_hd__decap_3 PHY_2108 ();
 sky130_fd_sc_hd__decap_3 PHY_2109 ();
 sky130_fd_sc_hd__decap_3 PHY_2110 ();
 sky130_fd_sc_hd__decap_3 PHY_2111 ();
 sky130_fd_sc_hd__decap_3 PHY_2112 ();
 sky130_fd_sc_hd__decap_3 PHY_2113 ();
 sky130_fd_sc_hd__decap_3 PHY_2114 ();
 sky130_fd_sc_hd__decap_3 PHY_2115 ();
 sky130_fd_sc_hd__decap_3 PHY_2116 ();
 sky130_fd_sc_hd__decap_3 PHY_2117 ();
 sky130_fd_sc_hd__decap_3 PHY_2118 ();
 sky130_fd_sc_hd__decap_3 PHY_2119 ();
 sky130_fd_sc_hd__decap_3 PHY_2120 ();
 sky130_fd_sc_hd__decap_3 PHY_2121 ();
 sky130_fd_sc_hd__decap_3 PHY_2122 ();
 sky130_fd_sc_hd__decap_3 PHY_2123 ();
 sky130_fd_sc_hd__decap_3 PHY_2124 ();
 sky130_fd_sc_hd__decap_3 PHY_2125 ();
 sky130_fd_sc_hd__decap_3 PHY_2126 ();
 sky130_fd_sc_hd__decap_3 PHY_2127 ();
 sky130_fd_sc_hd__decap_3 PHY_2128 ();
 sky130_fd_sc_hd__decap_3 PHY_2129 ();
 sky130_fd_sc_hd__decap_3 PHY_2130 ();
 sky130_fd_sc_hd__decap_3 PHY_2131 ();
 sky130_fd_sc_hd__decap_3 PHY_2132 ();
 sky130_fd_sc_hd__decap_3 PHY_2133 ();
 sky130_fd_sc_hd__decap_3 PHY_2134 ();
 sky130_fd_sc_hd__decap_3 PHY_2135 ();
 sky130_fd_sc_hd__decap_3 PHY_2136 ();
 sky130_fd_sc_hd__decap_3 PHY_2137 ();
 sky130_fd_sc_hd__decap_3 PHY_2138 ();
 sky130_fd_sc_hd__decap_3 PHY_2139 ();
 sky130_fd_sc_hd__decap_3 PHY_2140 ();
 sky130_fd_sc_hd__decap_3 PHY_2141 ();
 sky130_fd_sc_hd__decap_3 PHY_2142 ();
 sky130_fd_sc_hd__decap_3 PHY_2143 ();
 sky130_fd_sc_hd__decap_3 PHY_2144 ();
 sky130_fd_sc_hd__decap_3 PHY_2145 ();
 sky130_fd_sc_hd__decap_3 PHY_2146 ();
 sky130_fd_sc_hd__decap_3 PHY_2147 ();
 sky130_fd_sc_hd__decap_3 PHY_2148 ();
 sky130_fd_sc_hd__decap_3 PHY_2149 ();
 sky130_fd_sc_hd__decap_3 PHY_2150 ();
 sky130_fd_sc_hd__decap_3 PHY_2151 ();
 sky130_fd_sc_hd__decap_3 PHY_2152 ();
 sky130_fd_sc_hd__decap_3 PHY_2153 ();
 sky130_fd_sc_hd__decap_3 PHY_2154 ();
 sky130_fd_sc_hd__decap_3 PHY_2155 ();
 sky130_fd_sc_hd__decap_3 PHY_2156 ();
 sky130_fd_sc_hd__decap_3 PHY_2157 ();
 sky130_fd_sc_hd__decap_3 PHY_2158 ();
 sky130_fd_sc_hd__decap_3 PHY_2159 ();
 sky130_fd_sc_hd__decap_3 PHY_2160 ();
 sky130_fd_sc_hd__decap_3 PHY_2161 ();
 sky130_fd_sc_hd__decap_3 PHY_2162 ();
 sky130_fd_sc_hd__decap_3 PHY_2163 ();
 sky130_fd_sc_hd__decap_3 PHY_2164 ();
 sky130_fd_sc_hd__decap_3 PHY_2165 ();
 sky130_fd_sc_hd__decap_3 PHY_2166 ();
 sky130_fd_sc_hd__decap_3 PHY_2167 ();
 sky130_fd_sc_hd__decap_3 PHY_2168 ();
 sky130_fd_sc_hd__decap_3 PHY_2169 ();
 sky130_fd_sc_hd__decap_3 PHY_2170 ();
 sky130_fd_sc_hd__decap_3 PHY_2171 ();
 sky130_fd_sc_hd__decap_3 PHY_2172 ();
 sky130_fd_sc_hd__decap_3 PHY_2173 ();
 sky130_fd_sc_hd__decap_3 PHY_2174 ();
 sky130_fd_sc_hd__decap_3 PHY_2175 ();
 sky130_fd_sc_hd__decap_3 PHY_2176 ();
 sky130_fd_sc_hd__decap_3 PHY_2177 ();
 sky130_fd_sc_hd__decap_3 PHY_2178 ();
 sky130_fd_sc_hd__decap_3 PHY_2179 ();
 sky130_fd_sc_hd__decap_3 PHY_2180 ();
 sky130_fd_sc_hd__decap_3 PHY_2181 ();
 sky130_fd_sc_hd__decap_3 PHY_2182 ();
 sky130_fd_sc_hd__decap_3 PHY_2183 ();
 sky130_fd_sc_hd__decap_3 PHY_2184 ();
 sky130_fd_sc_hd__decap_3 PHY_2185 ();
 sky130_fd_sc_hd__decap_3 PHY_2186 ();
 sky130_fd_sc_hd__decap_3 PHY_2187 ();
 sky130_fd_sc_hd__decap_3 PHY_2188 ();
 sky130_fd_sc_hd__decap_3 PHY_2189 ();
 sky130_fd_sc_hd__decap_3 PHY_2190 ();
 sky130_fd_sc_hd__decap_3 PHY_2191 ();
 sky130_fd_sc_hd__decap_3 PHY_2192 ();
 sky130_fd_sc_hd__decap_3 PHY_2193 ();
 sky130_fd_sc_hd__decap_3 PHY_2194 ();
 sky130_fd_sc_hd__decap_3 PHY_2195 ();
 sky130_fd_sc_hd__decap_3 PHY_2196 ();
 sky130_fd_sc_hd__decap_3 PHY_2197 ();
 sky130_fd_sc_hd__decap_3 PHY_2198 ();
 sky130_fd_sc_hd__decap_3 PHY_2199 ();
 sky130_fd_sc_hd__decap_3 PHY_2200 ();
 sky130_fd_sc_hd__decap_3 PHY_2201 ();
 sky130_fd_sc_hd__decap_3 PHY_2202 ();
 sky130_fd_sc_hd__decap_3 PHY_2203 ();
 sky130_fd_sc_hd__decap_3 PHY_2204 ();
 sky130_fd_sc_hd__decap_3 PHY_2205 ();
 sky130_fd_sc_hd__decap_3 PHY_2206 ();
 sky130_fd_sc_hd__decap_3 PHY_2207 ();
 sky130_fd_sc_hd__decap_3 PHY_2208 ();
 sky130_fd_sc_hd__decap_3 PHY_2209 ();
 sky130_fd_sc_hd__decap_3 PHY_2210 ();
 sky130_fd_sc_hd__decap_3 PHY_2211 ();
 sky130_fd_sc_hd__decap_3 PHY_2212 ();
 sky130_fd_sc_hd__decap_3 PHY_2213 ();
 sky130_fd_sc_hd__decap_3 PHY_2214 ();
 sky130_fd_sc_hd__decap_3 PHY_2215 ();
 sky130_fd_sc_hd__decap_3 PHY_2216 ();
 sky130_fd_sc_hd__decap_3 PHY_2217 ();
 sky130_fd_sc_hd__decap_3 PHY_2218 ();
 sky130_fd_sc_hd__decap_3 PHY_2219 ();
 sky130_fd_sc_hd__decap_3 PHY_2220 ();
 sky130_fd_sc_hd__decap_3 PHY_2221 ();
 sky130_fd_sc_hd__decap_3 PHY_2222 ();
 sky130_fd_sc_hd__decap_3 PHY_2223 ();
 sky130_fd_sc_hd__decap_3 PHY_2224 ();
 sky130_fd_sc_hd__decap_3 PHY_2225 ();
 sky130_fd_sc_hd__decap_3 PHY_2226 ();
 sky130_fd_sc_hd__decap_3 PHY_2227 ();
 sky130_fd_sc_hd__decap_3 PHY_2228 ();
 sky130_fd_sc_hd__decap_3 PHY_2229 ();
 sky130_fd_sc_hd__decap_3 PHY_2230 ();
 sky130_fd_sc_hd__decap_3 PHY_2231 ();
 sky130_fd_sc_hd__decap_3 PHY_2232 ();
 sky130_fd_sc_hd__decap_3 PHY_2233 ();
 sky130_fd_sc_hd__decap_3 PHY_2234 ();
 sky130_fd_sc_hd__decap_3 PHY_2235 ();
 sky130_fd_sc_hd__decap_3 PHY_2236 ();
 sky130_fd_sc_hd__decap_3 PHY_2237 ();
 sky130_fd_sc_hd__decap_3 PHY_2238 ();
 sky130_fd_sc_hd__decap_3 PHY_2239 ();
 sky130_fd_sc_hd__decap_3 PHY_2240 ();
 sky130_fd_sc_hd__decap_3 PHY_2241 ();
 sky130_fd_sc_hd__decap_3 PHY_2242 ();
 sky130_fd_sc_hd__decap_3 PHY_2243 ();
 sky130_fd_sc_hd__decap_3 PHY_2244 ();
 sky130_fd_sc_hd__decap_3 PHY_2245 ();
 sky130_fd_sc_hd__decap_3 PHY_2246 ();
 sky130_fd_sc_hd__decap_3 PHY_2247 ();
 sky130_fd_sc_hd__decap_3 PHY_2248 ();
 sky130_fd_sc_hd__decap_3 PHY_2249 ();
 sky130_fd_sc_hd__decap_3 PHY_2250 ();
 sky130_fd_sc_hd__decap_3 PHY_2251 ();
 sky130_fd_sc_hd__decap_3 PHY_2252 ();
 sky130_fd_sc_hd__decap_3 PHY_2253 ();
 sky130_fd_sc_hd__decap_3 PHY_2254 ();
 sky130_fd_sc_hd__decap_3 PHY_2255 ();
 sky130_fd_sc_hd__decap_3 PHY_2256 ();
 sky130_fd_sc_hd__decap_3 PHY_2257 ();
 sky130_fd_sc_hd__decap_3 PHY_2258 ();
 sky130_fd_sc_hd__decap_3 PHY_2259 ();
 sky130_fd_sc_hd__decap_3 PHY_2260 ();
 sky130_fd_sc_hd__decap_3 PHY_2261 ();
 sky130_fd_sc_hd__decap_3 PHY_2262 ();
 sky130_fd_sc_hd__decap_3 PHY_2263 ();
 sky130_fd_sc_hd__decap_3 PHY_2264 ();
 sky130_fd_sc_hd__decap_3 PHY_2265 ();
 sky130_fd_sc_hd__decap_3 PHY_2266 ();
 sky130_fd_sc_hd__decap_3 PHY_2267 ();
 sky130_fd_sc_hd__decap_3 PHY_2268 ();
 sky130_fd_sc_hd__decap_3 PHY_2269 ();
 sky130_fd_sc_hd__decap_3 PHY_2270 ();
 sky130_fd_sc_hd__decap_3 PHY_2271 ();
 sky130_fd_sc_hd__decap_3 PHY_2272 ();
 sky130_fd_sc_hd__decap_3 PHY_2273 ();
 sky130_fd_sc_hd__decap_3 PHY_2274 ();
 sky130_fd_sc_hd__decap_3 PHY_2275 ();
 sky130_fd_sc_hd__decap_3 PHY_2276 ();
 sky130_fd_sc_hd__decap_3 PHY_2277 ();
 sky130_fd_sc_hd__decap_3 PHY_2278 ();
 sky130_fd_sc_hd__decap_3 PHY_2279 ();
 sky130_fd_sc_hd__decap_3 PHY_2280 ();
 sky130_fd_sc_hd__decap_3 PHY_2281 ();
 sky130_fd_sc_hd__decap_3 PHY_2282 ();
 sky130_fd_sc_hd__decap_3 PHY_2283 ();
 sky130_fd_sc_hd__decap_3 PHY_2284 ();
 sky130_fd_sc_hd__decap_3 PHY_2285 ();
 sky130_fd_sc_hd__decap_3 PHY_2286 ();
 sky130_fd_sc_hd__decap_3 PHY_2287 ();
 sky130_fd_sc_hd__decap_3 PHY_2288 ();
 sky130_fd_sc_hd__decap_3 PHY_2289 ();
 sky130_fd_sc_hd__decap_3 PHY_2290 ();
 sky130_fd_sc_hd__decap_3 PHY_2291 ();
 sky130_fd_sc_hd__decap_3 PHY_2292 ();
 sky130_fd_sc_hd__decap_3 PHY_2293 ();
 sky130_fd_sc_hd__decap_3 PHY_2294 ();
 sky130_fd_sc_hd__decap_3 PHY_2295 ();
 sky130_fd_sc_hd__decap_3 PHY_2296 ();
 sky130_fd_sc_hd__decap_3 PHY_2297 ();
 sky130_fd_sc_hd__decap_3 PHY_2298 ();
 sky130_fd_sc_hd__decap_3 PHY_2299 ();
 sky130_fd_sc_hd__decap_3 PHY_2300 ();
 sky130_fd_sc_hd__decap_3 PHY_2301 ();
 sky130_fd_sc_hd__decap_3 PHY_2302 ();
 sky130_fd_sc_hd__decap_3 PHY_2303 ();
 sky130_fd_sc_hd__decap_3 PHY_2304 ();
 sky130_fd_sc_hd__decap_3 PHY_2305 ();
 sky130_fd_sc_hd__decap_3 PHY_2306 ();
 sky130_fd_sc_hd__decap_3 PHY_2307 ();
 sky130_fd_sc_hd__decap_3 PHY_2308 ();
 sky130_fd_sc_hd__decap_3 PHY_2309 ();
 sky130_fd_sc_hd__decap_3 PHY_2310 ();
 sky130_fd_sc_hd__decap_3 PHY_2311 ();
 sky130_fd_sc_hd__decap_3 PHY_2312 ();
 sky130_fd_sc_hd__decap_3 PHY_2313 ();
 sky130_fd_sc_hd__decap_3 PHY_2314 ();
 sky130_fd_sc_hd__decap_3 PHY_2315 ();
 sky130_fd_sc_hd__decap_3 PHY_2316 ();
 sky130_fd_sc_hd__decap_3 PHY_2317 ();
 sky130_fd_sc_hd__decap_3 PHY_2318 ();
 sky130_fd_sc_hd__decap_3 PHY_2319 ();
 sky130_fd_sc_hd__decap_3 PHY_2320 ();
 sky130_fd_sc_hd__decap_3 PHY_2321 ();
 sky130_fd_sc_hd__decap_3 PHY_2322 ();
 sky130_fd_sc_hd__decap_3 PHY_2323 ();
 sky130_fd_sc_hd__decap_3 PHY_2324 ();
 sky130_fd_sc_hd__decap_3 PHY_2325 ();
 sky130_fd_sc_hd__decap_3 PHY_2326 ();
 sky130_fd_sc_hd__decap_3 PHY_2327 ();
 sky130_fd_sc_hd__decap_3 PHY_2328 ();
 sky130_fd_sc_hd__decap_3 PHY_2329 ();
 sky130_fd_sc_hd__decap_3 PHY_2330 ();
 sky130_fd_sc_hd__decap_3 PHY_2331 ();
 sky130_fd_sc_hd__decap_3 PHY_2332 ();
 sky130_fd_sc_hd__decap_3 PHY_2333 ();
 sky130_fd_sc_hd__decap_3 PHY_2334 ();
 sky130_fd_sc_hd__decap_3 PHY_2335 ();
 sky130_fd_sc_hd__decap_3 PHY_2336 ();
 sky130_fd_sc_hd__decap_3 PHY_2337 ();
 sky130_fd_sc_hd__decap_3 PHY_2338 ();
 sky130_fd_sc_hd__decap_3 PHY_2339 ();
 sky130_fd_sc_hd__decap_3 PHY_2340 ();
 sky130_fd_sc_hd__decap_3 PHY_2341 ();
 sky130_fd_sc_hd__decap_3 PHY_2342 ();
 sky130_fd_sc_hd__decap_3 PHY_2343 ();
 sky130_fd_sc_hd__decap_3 PHY_2344 ();
 sky130_fd_sc_hd__decap_3 PHY_2345 ();
 sky130_fd_sc_hd__decap_3 PHY_2346 ();
 sky130_fd_sc_hd__decap_3 PHY_2347 ();
 sky130_fd_sc_hd__decap_3 PHY_2348 ();
 sky130_fd_sc_hd__decap_3 PHY_2349 ();
 sky130_fd_sc_hd__decap_3 PHY_2350 ();
 sky130_fd_sc_hd__decap_3 PHY_2351 ();
 sky130_fd_sc_hd__decap_3 PHY_2352 ();
 sky130_fd_sc_hd__decap_3 PHY_2353 ();
 sky130_fd_sc_hd__decap_3 PHY_2354 ();
 sky130_fd_sc_hd__decap_3 PHY_2355 ();
 sky130_fd_sc_hd__decap_3 PHY_2356 ();
 sky130_fd_sc_hd__decap_3 PHY_2357 ();
 sky130_fd_sc_hd__decap_3 PHY_2358 ();
 sky130_fd_sc_hd__decap_3 PHY_2359 ();
 sky130_fd_sc_hd__decap_3 PHY_2360 ();
 sky130_fd_sc_hd__decap_3 PHY_2361 ();
 sky130_fd_sc_hd__decap_3 PHY_2362 ();
 sky130_fd_sc_hd__decap_3 PHY_2363 ();
 sky130_fd_sc_hd__decap_3 PHY_2364 ();
 sky130_fd_sc_hd__decap_3 PHY_2365 ();
 sky130_fd_sc_hd__decap_3 PHY_2366 ();
 sky130_fd_sc_hd__decap_3 PHY_2367 ();
 sky130_fd_sc_hd__decap_3 PHY_2368 ();
 sky130_fd_sc_hd__decap_3 PHY_2369 ();
 sky130_fd_sc_hd__decap_3 PHY_2370 ();
 sky130_fd_sc_hd__decap_3 PHY_2371 ();
 sky130_fd_sc_hd__decap_3 PHY_2372 ();
 sky130_fd_sc_hd__decap_3 PHY_2373 ();
 sky130_fd_sc_hd__decap_3 PHY_2374 ();
 sky130_fd_sc_hd__decap_3 PHY_2375 ();
 sky130_fd_sc_hd__decap_3 PHY_2376 ();
 sky130_fd_sc_hd__decap_3 PHY_2377 ();
 sky130_fd_sc_hd__decap_3 PHY_2378 ();
 sky130_fd_sc_hd__decap_3 PHY_2379 ();
 sky130_fd_sc_hd__decap_3 PHY_2380 ();
 sky130_fd_sc_hd__decap_3 PHY_2381 ();
 sky130_fd_sc_hd__decap_3 PHY_2382 ();
 sky130_fd_sc_hd__decap_3 PHY_2383 ();
 sky130_fd_sc_hd__decap_3 PHY_2384 ();
 sky130_fd_sc_hd__decap_3 PHY_2385 ();
 sky130_fd_sc_hd__decap_3 PHY_2386 ();
 sky130_fd_sc_hd__decap_3 PHY_2387 ();
 sky130_fd_sc_hd__decap_3 PHY_2388 ();
 sky130_fd_sc_hd__decap_3 PHY_2389 ();
 sky130_fd_sc_hd__decap_3 PHY_2390 ();
 sky130_fd_sc_hd__decap_3 PHY_2391 ();
 sky130_fd_sc_hd__decap_3 PHY_2392 ();
 sky130_fd_sc_hd__decap_3 PHY_2393 ();
 sky130_fd_sc_hd__decap_3 PHY_2394 ();
 sky130_fd_sc_hd__decap_3 PHY_2395 ();
 sky130_fd_sc_hd__decap_3 PHY_2396 ();
 sky130_fd_sc_hd__decap_3 PHY_2397 ();
 sky130_fd_sc_hd__decap_3 PHY_2398 ();
 sky130_fd_sc_hd__decap_3 PHY_2399 ();
 sky130_fd_sc_hd__decap_3 PHY_2400 ();
 sky130_fd_sc_hd__decap_3 PHY_2401 ();
 sky130_fd_sc_hd__decap_3 PHY_2402 ();
 sky130_fd_sc_hd__decap_3 PHY_2403 ();
 sky130_fd_sc_hd__decap_3 PHY_2404 ();
 sky130_fd_sc_hd__decap_3 PHY_2405 ();
 sky130_fd_sc_hd__decap_3 PHY_2406 ();
 sky130_fd_sc_hd__decap_3 PHY_2407 ();
 sky130_fd_sc_hd__decap_3 PHY_2408 ();
 sky130_fd_sc_hd__decap_3 PHY_2409 ();
 sky130_fd_sc_hd__decap_3 PHY_2410 ();
 sky130_fd_sc_hd__decap_3 PHY_2411 ();
 sky130_fd_sc_hd__decap_3 PHY_2412 ();
 sky130_fd_sc_hd__decap_3 PHY_2413 ();
 sky130_fd_sc_hd__decap_3 PHY_2414 ();
 sky130_fd_sc_hd__decap_3 PHY_2415 ();
 sky130_fd_sc_hd__decap_3 PHY_2416 ();
 sky130_fd_sc_hd__decap_3 PHY_2417 ();
 sky130_fd_sc_hd__decap_3 PHY_2418 ();
 sky130_fd_sc_hd__decap_3 PHY_2419 ();
 sky130_fd_sc_hd__decap_3 PHY_2420 ();
 sky130_fd_sc_hd__decap_3 PHY_2421 ();
 sky130_fd_sc_hd__decap_3 PHY_2422 ();
 sky130_fd_sc_hd__decap_3 PHY_2423 ();
 sky130_fd_sc_hd__decap_3 PHY_2424 ();
 sky130_fd_sc_hd__decap_3 PHY_2425 ();
 sky130_fd_sc_hd__decap_3 PHY_2426 ();
 sky130_fd_sc_hd__decap_3 PHY_2427 ();
 sky130_fd_sc_hd__decap_3 PHY_2428 ();
 sky130_fd_sc_hd__decap_3 PHY_2429 ();
 sky130_fd_sc_hd__decap_3 PHY_2430 ();
 sky130_fd_sc_hd__decap_3 PHY_2431 ();
 sky130_fd_sc_hd__decap_3 PHY_2432 ();
 sky130_fd_sc_hd__decap_3 PHY_2433 ();
 sky130_fd_sc_hd__decap_3 PHY_2434 ();
 sky130_fd_sc_hd__decap_3 PHY_2435 ();
 sky130_fd_sc_hd__decap_3 PHY_2436 ();
 sky130_fd_sc_hd__decap_3 PHY_2437 ();
 sky130_fd_sc_hd__decap_3 PHY_2438 ();
 sky130_fd_sc_hd__decap_3 PHY_2439 ();
 sky130_fd_sc_hd__decap_3 PHY_2440 ();
 sky130_fd_sc_hd__decap_3 PHY_2441 ();
 sky130_fd_sc_hd__decap_3 PHY_2442 ();
 sky130_fd_sc_hd__decap_3 PHY_2443 ();
 sky130_fd_sc_hd__decap_3 PHY_2444 ();
 sky130_fd_sc_hd__decap_3 PHY_2445 ();
 sky130_fd_sc_hd__decap_3 PHY_2446 ();
 sky130_fd_sc_hd__decap_3 PHY_2447 ();
 sky130_fd_sc_hd__decap_3 PHY_2448 ();
 sky130_fd_sc_hd__decap_3 PHY_2449 ();
 sky130_fd_sc_hd__decap_3 PHY_2450 ();
 sky130_fd_sc_hd__decap_3 PHY_2451 ();
 sky130_fd_sc_hd__decap_3 PHY_2452 ();
 sky130_fd_sc_hd__decap_3 PHY_2453 ();
 sky130_fd_sc_hd__decap_3 PHY_2454 ();
 sky130_fd_sc_hd__decap_3 PHY_2455 ();
 sky130_fd_sc_hd__decap_3 PHY_2456 ();
 sky130_fd_sc_hd__decap_3 PHY_2457 ();
 sky130_fd_sc_hd__decap_3 PHY_2458 ();
 sky130_fd_sc_hd__decap_3 PHY_2459 ();
 sky130_fd_sc_hd__decap_3 PHY_2460 ();
 sky130_fd_sc_hd__decap_3 PHY_2461 ();
 sky130_fd_sc_hd__decap_3 PHY_2462 ();
 sky130_fd_sc_hd__decap_3 PHY_2463 ();
 sky130_fd_sc_hd__decap_3 PHY_2464 ();
 sky130_fd_sc_hd__decap_3 PHY_2465 ();
 sky130_fd_sc_hd__decap_3 PHY_2466 ();
 sky130_fd_sc_hd__decap_3 PHY_2467 ();
 sky130_fd_sc_hd__decap_3 PHY_2468 ();
 sky130_fd_sc_hd__decap_3 PHY_2469 ();
 sky130_fd_sc_hd__decap_3 PHY_2470 ();
 sky130_fd_sc_hd__decap_3 PHY_2471 ();
 sky130_fd_sc_hd__decap_3 PHY_2472 ();
 sky130_fd_sc_hd__decap_3 PHY_2473 ();
 sky130_fd_sc_hd__decap_3 PHY_2474 ();
 sky130_fd_sc_hd__decap_3 PHY_2475 ();
 sky130_fd_sc_hd__decap_3 PHY_2476 ();
 sky130_fd_sc_hd__decap_3 PHY_2477 ();
 sky130_fd_sc_hd__decap_3 PHY_2478 ();
 sky130_fd_sc_hd__decap_3 PHY_2479 ();
 sky130_fd_sc_hd__decap_3 PHY_2480 ();
 sky130_fd_sc_hd__decap_3 PHY_2481 ();
 sky130_fd_sc_hd__decap_3 PHY_2482 ();
 sky130_fd_sc_hd__decap_3 PHY_2483 ();
 sky130_fd_sc_hd__decap_3 PHY_2484 ();
 sky130_fd_sc_hd__decap_3 PHY_2485 ();
 sky130_fd_sc_hd__decap_3 PHY_2486 ();
 sky130_fd_sc_hd__decap_3 PHY_2487 ();
 sky130_fd_sc_hd__decap_3 PHY_2488 ();
 sky130_fd_sc_hd__decap_3 PHY_2489 ();
 sky130_fd_sc_hd__decap_3 PHY_2490 ();
 sky130_fd_sc_hd__decap_3 PHY_2491 ();
 sky130_fd_sc_hd__decap_3 PHY_2492 ();
 sky130_fd_sc_hd__decap_3 PHY_2493 ();
 sky130_fd_sc_hd__decap_3 PHY_2494 ();
 sky130_fd_sc_hd__decap_3 PHY_2495 ();
 sky130_fd_sc_hd__decap_3 PHY_2496 ();
 sky130_fd_sc_hd__decap_3 PHY_2497 ();
 sky130_fd_sc_hd__decap_3 PHY_2498 ();
 sky130_fd_sc_hd__decap_3 PHY_2499 ();
 sky130_fd_sc_hd__decap_3 PHY_2500 ();
 sky130_fd_sc_hd__decap_3 PHY_2501 ();
 sky130_fd_sc_hd__decap_3 PHY_2502 ();
 sky130_fd_sc_hd__decap_3 PHY_2503 ();
 sky130_fd_sc_hd__decap_3 PHY_2504 ();
 sky130_fd_sc_hd__decap_3 PHY_2505 ();
 sky130_fd_sc_hd__decap_3 PHY_2506 ();
 sky130_fd_sc_hd__decap_3 PHY_2507 ();
 sky130_fd_sc_hd__decap_3 PHY_2508 ();
 sky130_fd_sc_hd__decap_3 PHY_2509 ();
 sky130_fd_sc_hd__decap_3 PHY_2510 ();
 sky130_fd_sc_hd__decap_3 PHY_2511 ();
 sky130_fd_sc_hd__decap_3 PHY_2512 ();
 sky130_fd_sc_hd__decap_3 PHY_2513 ();
 sky130_fd_sc_hd__decap_3 PHY_2514 ();
 sky130_fd_sc_hd__decap_3 PHY_2515 ();
 sky130_fd_sc_hd__decap_3 PHY_2516 ();
 sky130_fd_sc_hd__decap_3 PHY_2517 ();
 sky130_fd_sc_hd__decap_3 PHY_2518 ();
 sky130_fd_sc_hd__decap_3 PHY_2519 ();
 sky130_fd_sc_hd__decap_3 PHY_2520 ();
 sky130_fd_sc_hd__decap_3 PHY_2521 ();
 sky130_fd_sc_hd__decap_3 PHY_2522 ();
 sky130_fd_sc_hd__decap_3 PHY_2523 ();
 sky130_fd_sc_hd__decap_3 PHY_2524 ();
 sky130_fd_sc_hd__decap_3 PHY_2525 ();
 sky130_fd_sc_hd__decap_3 PHY_2526 ();
 sky130_fd_sc_hd__decap_3 PHY_2527 ();
 sky130_fd_sc_hd__decap_3 PHY_2528 ();
 sky130_fd_sc_hd__decap_3 PHY_2529 ();
 sky130_fd_sc_hd__decap_3 PHY_2530 ();
 sky130_fd_sc_hd__decap_3 PHY_2531 ();
 sky130_fd_sc_hd__decap_3 PHY_2532 ();
 sky130_fd_sc_hd__decap_3 PHY_2533 ();
 sky130_fd_sc_hd__decap_3 PHY_2534 ();
 sky130_fd_sc_hd__decap_3 PHY_2535 ();
 sky130_fd_sc_hd__decap_3 PHY_2536 ();
 sky130_fd_sc_hd__decap_3 PHY_2537 ();
 sky130_fd_sc_hd__decap_3 PHY_2538 ();
 sky130_fd_sc_hd__decap_3 PHY_2539 ();
 sky130_fd_sc_hd__decap_3 PHY_2540 ();
 sky130_fd_sc_hd__decap_3 PHY_2541 ();
 sky130_fd_sc_hd__decap_3 PHY_2542 ();
 sky130_fd_sc_hd__decap_3 PHY_2543 ();
 sky130_fd_sc_hd__decap_3 PHY_2544 ();
 sky130_fd_sc_hd__decap_3 PHY_2545 ();
 sky130_fd_sc_hd__decap_3 PHY_2546 ();
 sky130_fd_sc_hd__decap_3 PHY_2547 ();
 sky130_fd_sc_hd__decap_3 PHY_2548 ();
 sky130_fd_sc_hd__decap_3 PHY_2549 ();
 sky130_fd_sc_hd__decap_3 PHY_2550 ();
 sky130_fd_sc_hd__decap_3 PHY_2551 ();
 sky130_fd_sc_hd__decap_3 PHY_2552 ();
 sky130_fd_sc_hd__decap_3 PHY_2553 ();
 sky130_fd_sc_hd__decap_3 PHY_2554 ();
 sky130_fd_sc_hd__decap_3 PHY_2555 ();
 sky130_fd_sc_hd__decap_3 PHY_2556 ();
 sky130_fd_sc_hd__decap_3 PHY_2557 ();
 sky130_fd_sc_hd__decap_3 PHY_2558 ();
 sky130_fd_sc_hd__decap_3 PHY_2559 ();
 sky130_fd_sc_hd__decap_3 PHY_2560 ();
 sky130_fd_sc_hd__decap_3 PHY_2561 ();
 sky130_fd_sc_hd__decap_3 PHY_2562 ();
 sky130_fd_sc_hd__decap_3 PHY_2563 ();
 sky130_fd_sc_hd__decap_3 PHY_2564 ();
 sky130_fd_sc_hd__decap_3 PHY_2565 ();
 sky130_fd_sc_hd__decap_3 PHY_2566 ();
 sky130_fd_sc_hd__decap_3 PHY_2567 ();
 sky130_fd_sc_hd__decap_3 PHY_2568 ();
 sky130_fd_sc_hd__decap_3 PHY_2569 ();
 sky130_fd_sc_hd__decap_3 PHY_2570 ();
 sky130_fd_sc_hd__decap_3 PHY_2571 ();
 sky130_fd_sc_hd__decap_3 PHY_2572 ();
 sky130_fd_sc_hd__decap_3 PHY_2573 ();
 sky130_fd_sc_hd__decap_3 PHY_2574 ();
 sky130_fd_sc_hd__decap_3 PHY_2575 ();
 sky130_fd_sc_hd__decap_3 PHY_2576 ();
 sky130_fd_sc_hd__decap_3 PHY_2577 ();
 sky130_fd_sc_hd__decap_3 PHY_2578 ();
 sky130_fd_sc_hd__decap_3 PHY_2579 ();
 sky130_fd_sc_hd__decap_3 PHY_2580 ();
 sky130_fd_sc_hd__decap_3 PHY_2581 ();
 sky130_fd_sc_hd__decap_3 PHY_2582 ();
 sky130_fd_sc_hd__decap_3 PHY_2583 ();
 sky130_fd_sc_hd__decap_3 PHY_2584 ();
 sky130_fd_sc_hd__decap_3 PHY_2585 ();
 sky130_fd_sc_hd__decap_3 PHY_2586 ();
 sky130_fd_sc_hd__decap_3 PHY_2587 ();
 sky130_fd_sc_hd__decap_3 PHY_2588 ();
 sky130_fd_sc_hd__decap_3 PHY_2589 ();
 sky130_fd_sc_hd__decap_3 PHY_2590 ();
 sky130_fd_sc_hd__decap_3 PHY_2591 ();
 sky130_fd_sc_hd__decap_3 PHY_2592 ();
 sky130_fd_sc_hd__decap_3 PHY_2593 ();
 sky130_fd_sc_hd__decap_3 PHY_2594 ();
 sky130_fd_sc_hd__decap_3 PHY_2595 ();
 sky130_fd_sc_hd__decap_3 PHY_2596 ();
 sky130_fd_sc_hd__decap_3 PHY_2597 ();
 sky130_fd_sc_hd__decap_3 PHY_2598 ();
 sky130_fd_sc_hd__decap_3 PHY_2599 ();
 sky130_fd_sc_hd__decap_3 PHY_2600 ();
 sky130_fd_sc_hd__decap_3 PHY_2601 ();
 sky130_fd_sc_hd__decap_3 PHY_2602 ();
 sky130_fd_sc_hd__decap_3 PHY_2603 ();
 sky130_fd_sc_hd__decap_3 PHY_2604 ();
 sky130_fd_sc_hd__decap_3 PHY_2605 ();
 sky130_fd_sc_hd__decap_3 PHY_2606 ();
 sky130_fd_sc_hd__decap_3 PHY_2607 ();
 sky130_fd_sc_hd__decap_3 PHY_2608 ();
 sky130_fd_sc_hd__decap_3 PHY_2609 ();
 sky130_fd_sc_hd__decap_3 PHY_2610 ();
 sky130_fd_sc_hd__decap_3 PHY_2611 ();
 sky130_fd_sc_hd__decap_3 PHY_2612 ();
 sky130_fd_sc_hd__decap_3 PHY_2613 ();
 sky130_fd_sc_hd__decap_3 PHY_2614 ();
 sky130_fd_sc_hd__decap_3 PHY_2615 ();
 sky130_fd_sc_hd__decap_3 PHY_2616 ();
 sky130_fd_sc_hd__decap_3 PHY_2617 ();
 sky130_fd_sc_hd__decap_3 PHY_2618 ();
 sky130_fd_sc_hd__decap_3 PHY_2619 ();
 sky130_fd_sc_hd__decap_3 PHY_2620 ();
 sky130_fd_sc_hd__decap_3 PHY_2621 ();
 sky130_fd_sc_hd__decap_3 PHY_2622 ();
 sky130_fd_sc_hd__decap_3 PHY_2623 ();
 sky130_fd_sc_hd__decap_3 PHY_2624 ();
 sky130_fd_sc_hd__decap_3 PHY_2625 ();
 sky130_fd_sc_hd__decap_3 PHY_2626 ();
 sky130_fd_sc_hd__decap_3 PHY_2627 ();
 sky130_fd_sc_hd__decap_3 PHY_2628 ();
 sky130_fd_sc_hd__decap_3 PHY_2629 ();
 sky130_fd_sc_hd__decap_3 PHY_2630 ();
 sky130_fd_sc_hd__decap_3 PHY_2631 ();
 sky130_fd_sc_hd__decap_3 PHY_2632 ();
 sky130_fd_sc_hd__decap_3 PHY_2633 ();
 sky130_fd_sc_hd__decap_3 PHY_2634 ();
 sky130_fd_sc_hd__decap_3 PHY_2635 ();
 sky130_fd_sc_hd__decap_3 PHY_2636 ();
 sky130_fd_sc_hd__decap_3 PHY_2637 ();
 sky130_fd_sc_hd__decap_3 PHY_2638 ();
 sky130_fd_sc_hd__decap_3 PHY_2639 ();
 sky130_fd_sc_hd__decap_3 PHY_2640 ();
 sky130_fd_sc_hd__decap_3 PHY_2641 ();
 sky130_fd_sc_hd__decap_3 PHY_2642 ();
 sky130_fd_sc_hd__decap_3 PHY_2643 ();
 sky130_fd_sc_hd__decap_3 PHY_2644 ();
 sky130_fd_sc_hd__decap_3 PHY_2645 ();
 sky130_fd_sc_hd__decap_3 PHY_2646 ();
 sky130_fd_sc_hd__decap_3 PHY_2647 ();
 sky130_fd_sc_hd__decap_3 PHY_2648 ();
 sky130_fd_sc_hd__decap_3 PHY_2649 ();
 sky130_fd_sc_hd__decap_3 PHY_2650 ();
 sky130_fd_sc_hd__decap_3 PHY_2651 ();
 sky130_fd_sc_hd__decap_3 PHY_2652 ();
 sky130_fd_sc_hd__decap_3 PHY_2653 ();
 sky130_fd_sc_hd__decap_3 PHY_2654 ();
 sky130_fd_sc_hd__decap_3 PHY_2655 ();
 sky130_fd_sc_hd__decap_3 PHY_2656 ();
 sky130_fd_sc_hd__decap_3 PHY_2657 ();
 sky130_fd_sc_hd__decap_3 PHY_2658 ();
 sky130_fd_sc_hd__decap_3 PHY_2659 ();
 sky130_fd_sc_hd__decap_3 PHY_2660 ();
 sky130_fd_sc_hd__decap_3 PHY_2661 ();
 sky130_fd_sc_hd__decap_3 PHY_2662 ();
 sky130_fd_sc_hd__decap_3 PHY_2663 ();
 sky130_fd_sc_hd__decap_3 PHY_2664 ();
 sky130_fd_sc_hd__decap_3 PHY_2665 ();
 sky130_fd_sc_hd__decap_3 PHY_2666 ();
 sky130_fd_sc_hd__decap_3 PHY_2667 ();
 sky130_fd_sc_hd__decap_3 PHY_2668 ();
 sky130_fd_sc_hd__decap_3 PHY_2669 ();
 sky130_fd_sc_hd__decap_3 PHY_2670 ();
 sky130_fd_sc_hd__decap_3 PHY_2671 ();
 sky130_fd_sc_hd__decap_3 PHY_2672 ();
 sky130_fd_sc_hd__decap_3 PHY_2673 ();
 sky130_fd_sc_hd__decap_3 PHY_2674 ();
 sky130_fd_sc_hd__decap_3 PHY_2675 ();
 sky130_fd_sc_hd__decap_3 PHY_2676 ();
 sky130_fd_sc_hd__decap_3 PHY_2677 ();
 sky130_fd_sc_hd__decap_3 PHY_2678 ();
 sky130_fd_sc_hd__decap_3 PHY_2679 ();
 sky130_fd_sc_hd__decap_3 PHY_2680 ();
 sky130_fd_sc_hd__decap_3 PHY_2681 ();
 sky130_fd_sc_hd__decap_3 PHY_2682 ();
 sky130_fd_sc_hd__decap_3 PHY_2683 ();
 sky130_fd_sc_hd__decap_3 PHY_2684 ();
 sky130_fd_sc_hd__decap_3 PHY_2685 ();
 sky130_fd_sc_hd__decap_3 PHY_2686 ();
 sky130_fd_sc_hd__decap_3 PHY_2687 ();
 sky130_fd_sc_hd__decap_3 PHY_2688 ();
 sky130_fd_sc_hd__decap_3 PHY_2689 ();
 sky130_fd_sc_hd__decap_3 PHY_2690 ();
 sky130_fd_sc_hd__decap_3 PHY_2691 ();
 sky130_fd_sc_hd__decap_3 PHY_2692 ();
 sky130_fd_sc_hd__decap_3 PHY_2693 ();
 sky130_fd_sc_hd__decap_3 PHY_2694 ();
 sky130_fd_sc_hd__decap_3 PHY_2695 ();
 sky130_fd_sc_hd__decap_3 PHY_2696 ();
 sky130_fd_sc_hd__decap_3 PHY_2697 ();
 sky130_fd_sc_hd__decap_3 PHY_2698 ();
 sky130_fd_sc_hd__decap_3 PHY_2699 ();
 sky130_fd_sc_hd__decap_3 PHY_2700 ();
 sky130_fd_sc_hd__decap_3 PHY_2701 ();
 sky130_fd_sc_hd__decap_3 PHY_2702 ();
 sky130_fd_sc_hd__decap_3 PHY_2703 ();
 sky130_fd_sc_hd__decap_3 PHY_2704 ();
 sky130_fd_sc_hd__decap_3 PHY_2705 ();
 sky130_fd_sc_hd__decap_3 PHY_2706 ();
 sky130_fd_sc_hd__decap_3 PHY_2707 ();
 sky130_fd_sc_hd__decap_3 PHY_2708 ();
 sky130_fd_sc_hd__decap_3 PHY_2709 ();
 sky130_fd_sc_hd__decap_3 PHY_2710 ();
 sky130_fd_sc_hd__decap_3 PHY_2711 ();
 sky130_fd_sc_hd__decap_3 PHY_2712 ();
 sky130_fd_sc_hd__decap_3 PHY_2713 ();
 sky130_fd_sc_hd__decap_3 PHY_2714 ();
 sky130_fd_sc_hd__decap_3 PHY_2715 ();
 sky130_fd_sc_hd__decap_3 PHY_2716 ();
 sky130_fd_sc_hd__decap_3 PHY_2717 ();
 sky130_fd_sc_hd__decap_3 PHY_2718 ();
 sky130_fd_sc_hd__decap_3 PHY_2719 ();
 sky130_fd_sc_hd__decap_3 PHY_2720 ();
 sky130_fd_sc_hd__decap_3 PHY_2721 ();
 sky130_fd_sc_hd__decap_3 PHY_2722 ();
 sky130_fd_sc_hd__decap_3 PHY_2723 ();
 sky130_fd_sc_hd__decap_3 PHY_2724 ();
 sky130_fd_sc_hd__decap_3 PHY_2725 ();
 sky130_fd_sc_hd__decap_3 PHY_2726 ();
 sky130_fd_sc_hd__decap_3 PHY_2727 ();
 sky130_fd_sc_hd__decap_3 PHY_2728 ();
 sky130_fd_sc_hd__decap_3 PHY_2729 ();
 sky130_fd_sc_hd__decap_3 PHY_2730 ();
 sky130_fd_sc_hd__decap_3 PHY_2731 ();
 sky130_fd_sc_hd__decap_3 PHY_2732 ();
 sky130_fd_sc_hd__decap_3 PHY_2733 ();
 sky130_fd_sc_hd__decap_3 PHY_2734 ();
 sky130_fd_sc_hd__decap_3 PHY_2735 ();
 sky130_fd_sc_hd__decap_3 PHY_2736 ();
 sky130_fd_sc_hd__decap_3 PHY_2737 ();
 sky130_fd_sc_hd__decap_3 PHY_2738 ();
 sky130_fd_sc_hd__decap_3 PHY_2739 ();
 sky130_fd_sc_hd__decap_3 PHY_2740 ();
 sky130_fd_sc_hd__decap_3 PHY_2741 ();
 sky130_fd_sc_hd__decap_3 PHY_2742 ();
 sky130_fd_sc_hd__decap_3 PHY_2743 ();
 sky130_fd_sc_hd__decap_3 PHY_2744 ();
 sky130_fd_sc_hd__decap_3 PHY_2745 ();
 sky130_fd_sc_hd__decap_3 PHY_2746 ();
 sky130_fd_sc_hd__decap_3 PHY_2747 ();
 sky130_fd_sc_hd__decap_3 PHY_2748 ();
 sky130_fd_sc_hd__decap_3 PHY_2749 ();
 sky130_fd_sc_hd__decap_3 PHY_2750 ();
 sky130_fd_sc_hd__decap_3 PHY_2751 ();
 sky130_fd_sc_hd__decap_3 PHY_2752 ();
 sky130_fd_sc_hd__decap_3 PHY_2753 ();
 sky130_fd_sc_hd__decap_3 PHY_2754 ();
 sky130_fd_sc_hd__decap_3 PHY_2755 ();
 sky130_fd_sc_hd__decap_3 PHY_2756 ();
 sky130_fd_sc_hd__decap_3 PHY_2757 ();
 sky130_fd_sc_hd__decap_3 PHY_2758 ();
 sky130_fd_sc_hd__decap_3 PHY_2759 ();
 sky130_fd_sc_hd__decap_3 PHY_2760 ();
 sky130_fd_sc_hd__decap_3 PHY_2761 ();
 sky130_fd_sc_hd__decap_3 PHY_2762 ();
 sky130_fd_sc_hd__decap_3 PHY_2763 ();
 sky130_fd_sc_hd__decap_3 PHY_2764 ();
 sky130_fd_sc_hd__decap_3 PHY_2765 ();
 sky130_fd_sc_hd__decap_3 PHY_2766 ();
 sky130_fd_sc_hd__decap_3 PHY_2767 ();
 sky130_fd_sc_hd__decap_3 PHY_2768 ();
 sky130_fd_sc_hd__decap_3 PHY_2769 ();
 sky130_fd_sc_hd__decap_3 PHY_2770 ();
 sky130_fd_sc_hd__decap_3 PHY_2771 ();
 sky130_fd_sc_hd__decap_3 PHY_2772 ();
 sky130_fd_sc_hd__decap_3 PHY_2773 ();
 sky130_fd_sc_hd__decap_3 PHY_2774 ();
 sky130_fd_sc_hd__decap_3 PHY_2775 ();
 sky130_fd_sc_hd__decap_3 PHY_2776 ();
 sky130_fd_sc_hd__decap_3 PHY_2777 ();
 sky130_fd_sc_hd__decap_3 PHY_2778 ();
 sky130_fd_sc_hd__decap_3 PHY_2779 ();
 sky130_fd_sc_hd__decap_3 PHY_2780 ();
 sky130_fd_sc_hd__decap_3 PHY_2781 ();
 sky130_fd_sc_hd__decap_3 PHY_2782 ();
 sky130_fd_sc_hd__decap_3 PHY_2783 ();
 sky130_fd_sc_hd__decap_3 PHY_2784 ();
 sky130_fd_sc_hd__decap_3 PHY_2785 ();
 sky130_fd_sc_hd__decap_3 PHY_2786 ();
 sky130_fd_sc_hd__decap_3 PHY_2787 ();
 sky130_fd_sc_hd__decap_3 PHY_2788 ();
 sky130_fd_sc_hd__decap_3 PHY_2789 ();
 sky130_fd_sc_hd__decap_3 PHY_2790 ();
 sky130_fd_sc_hd__decap_3 PHY_2791 ();
 sky130_fd_sc_hd__decap_3 PHY_2792 ();
 sky130_fd_sc_hd__decap_3 PHY_2793 ();
 sky130_fd_sc_hd__decap_3 PHY_2794 ();
 sky130_fd_sc_hd__decap_3 PHY_2795 ();
 sky130_fd_sc_hd__decap_3 PHY_2796 ();
 sky130_fd_sc_hd__decap_3 PHY_2797 ();
 sky130_fd_sc_hd__decap_3 PHY_2798 ();
 sky130_fd_sc_hd__decap_3 PHY_2799 ();
 sky130_fd_sc_hd__decap_3 PHY_2800 ();
 sky130_fd_sc_hd__decap_3 PHY_2801 ();
 sky130_fd_sc_hd__decap_3 PHY_2802 ();
 sky130_fd_sc_hd__decap_3 PHY_2803 ();
 sky130_fd_sc_hd__decap_3 PHY_2804 ();
 sky130_fd_sc_hd__decap_3 PHY_2805 ();
 sky130_fd_sc_hd__decap_3 PHY_2806 ();
 sky130_fd_sc_hd__decap_3 PHY_2807 ();
 sky130_fd_sc_hd__decap_3 PHY_2808 ();
 sky130_fd_sc_hd__decap_3 PHY_2809 ();
 sky130_fd_sc_hd__decap_3 PHY_2810 ();
 sky130_fd_sc_hd__decap_3 PHY_2811 ();
 sky130_fd_sc_hd__decap_3 PHY_2812 ();
 sky130_fd_sc_hd__decap_3 PHY_2813 ();
 sky130_fd_sc_hd__decap_3 PHY_2814 ();
 sky130_fd_sc_hd__decap_3 PHY_2815 ();
 sky130_fd_sc_hd__decap_3 PHY_2816 ();
 sky130_fd_sc_hd__decap_3 PHY_2817 ();
 sky130_fd_sc_hd__decap_3 PHY_2818 ();
 sky130_fd_sc_hd__decap_3 PHY_2819 ();
 sky130_fd_sc_hd__decap_3 PHY_2820 ();
 sky130_fd_sc_hd__decap_3 PHY_2821 ();
 sky130_fd_sc_hd__decap_3 PHY_2822 ();
 sky130_fd_sc_hd__decap_3 PHY_2823 ();
 sky130_fd_sc_hd__decap_3 PHY_2824 ();
 sky130_fd_sc_hd__decap_3 PHY_2825 ();
 sky130_fd_sc_hd__decap_3 PHY_2826 ();
 sky130_fd_sc_hd__decap_3 PHY_2827 ();
 sky130_fd_sc_hd__decap_3 PHY_2828 ();
 sky130_fd_sc_hd__decap_3 PHY_2829 ();
 sky130_fd_sc_hd__decap_3 PHY_2830 ();
 sky130_fd_sc_hd__decap_3 PHY_2831 ();
 sky130_fd_sc_hd__decap_3 PHY_2832 ();
 sky130_fd_sc_hd__decap_3 PHY_2833 ();
 sky130_fd_sc_hd__decap_3 PHY_2834 ();
 sky130_fd_sc_hd__decap_3 PHY_2835 ();
 sky130_fd_sc_hd__decap_3 PHY_2836 ();
 sky130_fd_sc_hd__decap_3 PHY_2837 ();
 sky130_fd_sc_hd__decap_3 PHY_2838 ();
 sky130_fd_sc_hd__decap_3 PHY_2839 ();
 sky130_fd_sc_hd__decap_3 PHY_2840 ();
 sky130_fd_sc_hd__decap_3 PHY_2841 ();
 sky130_fd_sc_hd__decap_3 PHY_2842 ();
 sky130_fd_sc_hd__decap_3 PHY_2843 ();
 sky130_fd_sc_hd__decap_3 PHY_2844 ();
 sky130_fd_sc_hd__decap_3 PHY_2845 ();
 sky130_fd_sc_hd__decap_3 PHY_2846 ();
 sky130_fd_sc_hd__decap_3 PHY_2847 ();
 sky130_fd_sc_hd__decap_3 PHY_2848 ();
 sky130_fd_sc_hd__decap_3 PHY_2849 ();
 sky130_fd_sc_hd__decap_3 PHY_2850 ();
 sky130_fd_sc_hd__decap_3 PHY_2851 ();
 sky130_fd_sc_hd__decap_3 PHY_2852 ();
 sky130_fd_sc_hd__decap_3 PHY_2853 ();
 sky130_fd_sc_hd__decap_3 PHY_2854 ();
 sky130_fd_sc_hd__decap_3 PHY_2855 ();
 sky130_fd_sc_hd__decap_3 PHY_2856 ();
 sky130_fd_sc_hd__decap_3 PHY_2857 ();
 sky130_fd_sc_hd__decap_3 PHY_2858 ();
 sky130_fd_sc_hd__decap_3 PHY_2859 ();
 sky130_fd_sc_hd__decap_3 PHY_2860 ();
 sky130_fd_sc_hd__decap_3 PHY_2861 ();
 sky130_fd_sc_hd__decap_3 PHY_2862 ();
 sky130_fd_sc_hd__decap_3 PHY_2863 ();
 sky130_fd_sc_hd__decap_3 PHY_2864 ();
 sky130_fd_sc_hd__decap_3 PHY_2865 ();
 sky130_fd_sc_hd__decap_3 PHY_2866 ();
 sky130_fd_sc_hd__decap_3 PHY_2867 ();
 sky130_fd_sc_hd__decap_3 PHY_2868 ();
 sky130_fd_sc_hd__decap_3 PHY_2869 ();
 sky130_fd_sc_hd__decap_3 PHY_2870 ();
 sky130_fd_sc_hd__decap_3 PHY_2871 ();
 sky130_fd_sc_hd__decap_3 PHY_2872 ();
 sky130_fd_sc_hd__decap_3 PHY_2873 ();
 sky130_fd_sc_hd__decap_3 PHY_2874 ();
 sky130_fd_sc_hd__decap_3 PHY_2875 ();
 sky130_fd_sc_hd__decap_3 PHY_2876 ();
 sky130_fd_sc_hd__decap_3 PHY_2877 ();
 sky130_fd_sc_hd__decap_3 PHY_2878 ();
 sky130_fd_sc_hd__decap_3 PHY_2879 ();
 sky130_fd_sc_hd__decap_3 PHY_2880 ();
 sky130_fd_sc_hd__decap_3 PHY_2881 ();
 sky130_fd_sc_hd__decap_3 PHY_2882 ();
 sky130_fd_sc_hd__decap_3 PHY_2883 ();
 sky130_fd_sc_hd__decap_3 PHY_2884 ();
 sky130_fd_sc_hd__decap_3 PHY_2885 ();
 sky130_fd_sc_hd__decap_3 PHY_2886 ();
 sky130_fd_sc_hd__decap_3 PHY_2887 ();
 sky130_fd_sc_hd__decap_3 PHY_2888 ();
 sky130_fd_sc_hd__decap_3 PHY_2889 ();
 sky130_fd_sc_hd__decap_3 PHY_2890 ();
 sky130_fd_sc_hd__decap_3 PHY_2891 ();
 sky130_fd_sc_hd__decap_3 PHY_2892 ();
 sky130_fd_sc_hd__decap_3 PHY_2893 ();
 sky130_fd_sc_hd__decap_3 PHY_2894 ();
 sky130_fd_sc_hd__decap_3 PHY_2895 ();
 sky130_fd_sc_hd__decap_3 PHY_2896 ();
 sky130_fd_sc_hd__decap_3 PHY_2897 ();
 sky130_fd_sc_hd__decap_3 PHY_2898 ();
 sky130_fd_sc_hd__decap_3 PHY_2899 ();
 sky130_fd_sc_hd__decap_3 PHY_2900 ();
 sky130_fd_sc_hd__decap_3 PHY_2901 ();
 sky130_fd_sc_hd__decap_3 PHY_2902 ();
 sky130_fd_sc_hd__decap_3 PHY_2903 ();
 sky130_fd_sc_hd__decap_3 PHY_2904 ();
 sky130_fd_sc_hd__decap_3 PHY_2905 ();
 sky130_fd_sc_hd__decap_3 PHY_2906 ();
 sky130_fd_sc_hd__decap_3 PHY_2907 ();
 sky130_fd_sc_hd__decap_3 PHY_2908 ();
 sky130_fd_sc_hd__decap_3 PHY_2909 ();
 sky130_fd_sc_hd__decap_3 PHY_2910 ();
 sky130_fd_sc_hd__decap_3 PHY_2911 ();
 sky130_fd_sc_hd__decap_3 PHY_2912 ();
 sky130_fd_sc_hd__decap_3 PHY_2913 ();
 sky130_fd_sc_hd__decap_3 PHY_2914 ();
 sky130_fd_sc_hd__decap_3 PHY_2915 ();
 sky130_fd_sc_hd__decap_3 PHY_2916 ();
 sky130_fd_sc_hd__decap_3 PHY_2917 ();
 sky130_fd_sc_hd__decap_3 PHY_2918 ();
 sky130_fd_sc_hd__decap_3 PHY_2919 ();
 sky130_fd_sc_hd__decap_3 PHY_2920 ();
 sky130_fd_sc_hd__decap_3 PHY_2921 ();
 sky130_fd_sc_hd__decap_3 PHY_2922 ();
 sky130_fd_sc_hd__decap_3 PHY_2923 ();
 sky130_fd_sc_hd__decap_3 PHY_2924 ();
 sky130_fd_sc_hd__decap_3 PHY_2925 ();
 sky130_fd_sc_hd__decap_3 PHY_2926 ();
 sky130_fd_sc_hd__decap_3 PHY_2927 ();
 sky130_fd_sc_hd__decap_3 PHY_2928 ();
 sky130_fd_sc_hd__decap_3 PHY_2929 ();
 sky130_fd_sc_hd__decap_3 PHY_2930 ();
 sky130_fd_sc_hd__decap_3 PHY_2931 ();
 sky130_fd_sc_hd__decap_3 PHY_2932 ();
 sky130_fd_sc_hd__decap_3 PHY_2933 ();
 sky130_fd_sc_hd__decap_3 PHY_2934 ();
 sky130_fd_sc_hd__decap_3 PHY_2935 ();
 sky130_fd_sc_hd__decap_3 PHY_2936 ();
 sky130_fd_sc_hd__decap_3 PHY_2937 ();
 sky130_fd_sc_hd__decap_3 PHY_2938 ();
 sky130_fd_sc_hd__decap_3 PHY_2939 ();
 sky130_fd_sc_hd__decap_3 PHY_2940 ();
 sky130_fd_sc_hd__decap_3 PHY_2941 ();
 sky130_fd_sc_hd__decap_3 PHY_2942 ();
 sky130_fd_sc_hd__decap_3 PHY_2943 ();
 sky130_fd_sc_hd__decap_3 PHY_2944 ();
 sky130_fd_sc_hd__decap_3 PHY_2945 ();
 sky130_fd_sc_hd__decap_3 PHY_2946 ();
 sky130_fd_sc_hd__decap_3 PHY_2947 ();
 sky130_fd_sc_hd__decap_3 PHY_2948 ();
 sky130_fd_sc_hd__decap_3 PHY_2949 ();
 sky130_fd_sc_hd__decap_3 PHY_2950 ();
 sky130_fd_sc_hd__decap_3 PHY_2951 ();
 sky130_fd_sc_hd__decap_3 PHY_2952 ();
 sky130_fd_sc_hd__decap_3 PHY_2953 ();
 sky130_fd_sc_hd__decap_3 PHY_2954 ();
 sky130_fd_sc_hd__decap_3 PHY_2955 ();
 sky130_fd_sc_hd__decap_3 PHY_2956 ();
 sky130_fd_sc_hd__decap_3 PHY_2957 ();
 sky130_fd_sc_hd__decap_3 PHY_2958 ();
 sky130_fd_sc_hd__decap_3 PHY_2959 ();
 sky130_fd_sc_hd__decap_3 PHY_2960 ();
 sky130_fd_sc_hd__decap_3 PHY_2961 ();
 sky130_fd_sc_hd__decap_3 PHY_2962 ();
 sky130_fd_sc_hd__decap_3 PHY_2963 ();
 sky130_fd_sc_hd__decap_3 PHY_2964 ();
 sky130_fd_sc_hd__decap_3 PHY_2965 ();
 sky130_fd_sc_hd__decap_3 PHY_2966 ();
 sky130_fd_sc_hd__decap_3 PHY_2967 ();
 sky130_fd_sc_hd__decap_3 PHY_2968 ();
 sky130_fd_sc_hd__decap_3 PHY_2969 ();
 sky130_fd_sc_hd__decap_3 PHY_2970 ();
 sky130_fd_sc_hd__decap_3 PHY_2971 ();
 sky130_fd_sc_hd__decap_3 PHY_2972 ();
 sky130_fd_sc_hd__decap_3 PHY_2973 ();
 sky130_fd_sc_hd__decap_3 PHY_2974 ();
 sky130_fd_sc_hd__decap_3 PHY_2975 ();
 sky130_fd_sc_hd__decap_3 PHY_2976 ();
 sky130_fd_sc_hd__decap_3 PHY_2977 ();
 sky130_fd_sc_hd__decap_3 PHY_2978 ();
 sky130_fd_sc_hd__decap_3 PHY_2979 ();
 sky130_fd_sc_hd__decap_3 PHY_2980 ();
 sky130_fd_sc_hd__decap_3 PHY_2981 ();
 sky130_fd_sc_hd__decap_3 PHY_2982 ();
 sky130_fd_sc_hd__decap_3 PHY_2983 ();
 sky130_fd_sc_hd__decap_3 PHY_2984 ();
 sky130_fd_sc_hd__decap_3 PHY_2985 ();
 sky130_fd_sc_hd__decap_3 PHY_2986 ();
 sky130_fd_sc_hd__decap_3 PHY_2987 ();
 sky130_fd_sc_hd__decap_3 PHY_2988 ();
 sky130_fd_sc_hd__decap_3 PHY_2989 ();
 sky130_fd_sc_hd__decap_3 PHY_2990 ();
 sky130_fd_sc_hd__decap_3 PHY_2991 ();
 sky130_fd_sc_hd__decap_3 PHY_2992 ();
 sky130_fd_sc_hd__decap_3 PHY_2993 ();
 sky130_fd_sc_hd__decap_3 PHY_2994 ();
 sky130_fd_sc_hd__decap_3 PHY_2995 ();
 sky130_fd_sc_hd__decap_3 PHY_2996 ();
 sky130_fd_sc_hd__decap_3 PHY_2997 ();
 sky130_fd_sc_hd__decap_3 PHY_2998 ();
 sky130_fd_sc_hd__decap_3 PHY_2999 ();
 sky130_fd_sc_hd__decap_3 PHY_3000 ();
 sky130_fd_sc_hd__decap_3 PHY_3001 ();
 sky130_fd_sc_hd__decap_3 PHY_3002 ();
 sky130_fd_sc_hd__decap_3 PHY_3003 ();
 sky130_fd_sc_hd__decap_3 PHY_3004 ();
 sky130_fd_sc_hd__decap_3 PHY_3005 ();
 sky130_fd_sc_hd__decap_3 PHY_3006 ();
 sky130_fd_sc_hd__decap_3 PHY_3007 ();
 sky130_fd_sc_hd__decap_3 PHY_3008 ();
 sky130_fd_sc_hd__decap_3 PHY_3009 ();
 sky130_fd_sc_hd__decap_3 PHY_3010 ();
 sky130_fd_sc_hd__decap_3 PHY_3011 ();
 sky130_fd_sc_hd__decap_3 PHY_3012 ();
 sky130_fd_sc_hd__decap_3 PHY_3013 ();
 sky130_fd_sc_hd__decap_3 PHY_3014 ();
 sky130_fd_sc_hd__decap_3 PHY_3015 ();
 sky130_fd_sc_hd__decap_3 PHY_3016 ();
 sky130_fd_sc_hd__decap_3 PHY_3017 ();
 sky130_fd_sc_hd__decap_3 PHY_3018 ();
 sky130_fd_sc_hd__decap_3 PHY_3019 ();
 sky130_fd_sc_hd__decap_3 PHY_3020 ();
 sky130_fd_sc_hd__decap_3 PHY_3021 ();
 sky130_fd_sc_hd__decap_3 PHY_3022 ();
 sky130_fd_sc_hd__decap_3 PHY_3023 ();
 sky130_fd_sc_hd__decap_3 PHY_3024 ();
 sky130_fd_sc_hd__decap_3 PHY_3025 ();
 sky130_fd_sc_hd__decap_3 PHY_3026 ();
 sky130_fd_sc_hd__decap_3 PHY_3027 ();
 sky130_fd_sc_hd__decap_3 PHY_3028 ();
 sky130_fd_sc_hd__decap_3 PHY_3029 ();
 sky130_fd_sc_hd__decap_3 PHY_3030 ();
 sky130_fd_sc_hd__decap_3 PHY_3031 ();
 sky130_fd_sc_hd__decap_3 PHY_3032 ();
 sky130_fd_sc_hd__decap_3 PHY_3033 ();
 sky130_fd_sc_hd__decap_3 PHY_3034 ();
 sky130_fd_sc_hd__decap_3 PHY_3035 ();
 sky130_fd_sc_hd__decap_3 PHY_3036 ();
 sky130_fd_sc_hd__decap_3 PHY_3037 ();
 sky130_fd_sc_hd__decap_3 PHY_3038 ();
 sky130_fd_sc_hd__decap_3 PHY_3039 ();
 sky130_fd_sc_hd__decap_3 PHY_3040 ();
 sky130_fd_sc_hd__decap_3 PHY_3041 ();
 sky130_fd_sc_hd__decap_3 PHY_3042 ();
 sky130_fd_sc_hd__decap_3 PHY_3043 ();
 sky130_fd_sc_hd__decap_3 PHY_3044 ();
 sky130_fd_sc_hd__decap_3 PHY_3045 ();
 sky130_fd_sc_hd__decap_3 PHY_3046 ();
 sky130_fd_sc_hd__decap_3 PHY_3047 ();
 sky130_fd_sc_hd__decap_3 PHY_3048 ();
 sky130_fd_sc_hd__decap_3 PHY_3049 ();
 sky130_fd_sc_hd__decap_3 PHY_3050 ();
 sky130_fd_sc_hd__decap_3 PHY_3051 ();
 sky130_fd_sc_hd__decap_3 PHY_3052 ();
 sky130_fd_sc_hd__decap_3 PHY_3053 ();
 sky130_fd_sc_hd__decap_3 PHY_3054 ();
 sky130_fd_sc_hd__decap_3 PHY_3055 ();
 sky130_fd_sc_hd__decap_3 PHY_3056 ();
 sky130_fd_sc_hd__decap_3 PHY_3057 ();
 sky130_fd_sc_hd__decap_3 PHY_3058 ();
 sky130_fd_sc_hd__decap_3 PHY_3059 ();
 sky130_fd_sc_hd__decap_3 PHY_3060 ();
 sky130_fd_sc_hd__decap_3 PHY_3061 ();
 sky130_fd_sc_hd__decap_3 PHY_3062 ();
 sky130_fd_sc_hd__decap_3 PHY_3063 ();
 sky130_fd_sc_hd__decap_3 PHY_3064 ();
 sky130_fd_sc_hd__decap_3 PHY_3065 ();
 sky130_fd_sc_hd__decap_3 PHY_3066 ();
 sky130_fd_sc_hd__decap_3 PHY_3067 ();
 sky130_fd_sc_hd__decap_3 PHY_3068 ();
 sky130_fd_sc_hd__decap_3 PHY_3069 ();
 sky130_fd_sc_hd__decap_3 PHY_3070 ();
 sky130_fd_sc_hd__decap_3 PHY_3071 ();
 sky130_fd_sc_hd__decap_3 PHY_3072 ();
 sky130_fd_sc_hd__decap_3 PHY_3073 ();
 sky130_fd_sc_hd__decap_3 PHY_3074 ();
 sky130_fd_sc_hd__decap_3 PHY_3075 ();
 sky130_fd_sc_hd__decap_3 PHY_3076 ();
 sky130_fd_sc_hd__decap_3 PHY_3077 ();
 sky130_fd_sc_hd__decap_3 PHY_3078 ();
 sky130_fd_sc_hd__decap_3 PHY_3079 ();
 sky130_fd_sc_hd__decap_3 PHY_3080 ();
 sky130_fd_sc_hd__decap_3 PHY_3081 ();
 sky130_fd_sc_hd__decap_3 PHY_3082 ();
 sky130_fd_sc_hd__decap_3 PHY_3083 ();
 sky130_fd_sc_hd__decap_3 PHY_3084 ();
 sky130_fd_sc_hd__decap_3 PHY_3085 ();
 sky130_fd_sc_hd__decap_3 PHY_3086 ();
 sky130_fd_sc_hd__decap_3 PHY_3087 ();
 sky130_fd_sc_hd__decap_3 PHY_3088 ();
 sky130_fd_sc_hd__decap_3 PHY_3089 ();
 sky130_fd_sc_hd__decap_3 PHY_3090 ();
 sky130_fd_sc_hd__decap_3 PHY_3091 ();
 sky130_fd_sc_hd__decap_3 PHY_3092 ();
 sky130_fd_sc_hd__decap_3 PHY_3093 ();
 sky130_fd_sc_hd__decap_3 PHY_3094 ();
 sky130_fd_sc_hd__decap_3 PHY_3095 ();
 sky130_fd_sc_hd__decap_3 PHY_3096 ();
 sky130_fd_sc_hd__decap_3 PHY_3097 ();
 sky130_fd_sc_hd__decap_3 PHY_3098 ();
 sky130_fd_sc_hd__decap_3 PHY_3099 ();
 sky130_fd_sc_hd__decap_3 PHY_3100 ();
 sky130_fd_sc_hd__decap_3 PHY_3101 ();
 sky130_fd_sc_hd__decap_3 PHY_3102 ();
 sky130_fd_sc_hd__decap_3 PHY_3103 ();
 sky130_fd_sc_hd__decap_3 PHY_3104 ();
 sky130_fd_sc_hd__decap_3 PHY_3105 ();
 sky130_fd_sc_hd__decap_3 PHY_3106 ();
 sky130_fd_sc_hd__decap_3 PHY_3107 ();
 sky130_fd_sc_hd__decap_3 PHY_3108 ();
 sky130_fd_sc_hd__decap_3 PHY_3109 ();
 sky130_fd_sc_hd__decap_3 PHY_3110 ();
 sky130_fd_sc_hd__decap_3 PHY_3111 ();
 sky130_fd_sc_hd__decap_3 PHY_3112 ();
 sky130_fd_sc_hd__decap_3 PHY_3113 ();
 sky130_fd_sc_hd__decap_3 PHY_3114 ();
 sky130_fd_sc_hd__decap_3 PHY_3115 ();
 sky130_fd_sc_hd__decap_3 PHY_3116 ();
 sky130_fd_sc_hd__decap_3 PHY_3117 ();
 sky130_fd_sc_hd__decap_3 PHY_3118 ();
 sky130_fd_sc_hd__decap_3 PHY_3119 ();
 sky130_fd_sc_hd__decap_3 PHY_3120 ();
 sky130_fd_sc_hd__decap_3 PHY_3121 ();
 sky130_fd_sc_hd__decap_3 PHY_3122 ();
 sky130_fd_sc_hd__decap_3 PHY_3123 ();
 sky130_fd_sc_hd__decap_3 PHY_3124 ();
 sky130_fd_sc_hd__decap_3 PHY_3125 ();
 sky130_fd_sc_hd__decap_3 PHY_3126 ();
 sky130_fd_sc_hd__decap_3 PHY_3127 ();
 sky130_fd_sc_hd__decap_3 PHY_3128 ();
 sky130_fd_sc_hd__decap_3 PHY_3129 ();
 sky130_fd_sc_hd__decap_3 PHY_3130 ();
 sky130_fd_sc_hd__decap_3 PHY_3131 ();
 sky130_fd_sc_hd__decap_3 PHY_3132 ();
 sky130_fd_sc_hd__decap_3 PHY_3133 ();
 sky130_fd_sc_hd__decap_3 PHY_3134 ();
 sky130_fd_sc_hd__decap_3 PHY_3135 ();
 sky130_fd_sc_hd__decap_3 PHY_3136 ();
 sky130_fd_sc_hd__decap_3 PHY_3137 ();
 sky130_fd_sc_hd__decap_3 PHY_3138 ();
 sky130_fd_sc_hd__decap_3 PHY_3139 ();
 sky130_fd_sc_hd__decap_3 PHY_3140 ();
 sky130_fd_sc_hd__decap_3 PHY_3141 ();
 sky130_fd_sc_hd__decap_3 PHY_3142 ();
 sky130_fd_sc_hd__decap_3 PHY_3143 ();
 sky130_fd_sc_hd__decap_3 PHY_3144 ();
 sky130_fd_sc_hd__decap_3 PHY_3145 ();
 sky130_fd_sc_hd__decap_3 PHY_3146 ();
 sky130_fd_sc_hd__decap_3 PHY_3147 ();
 sky130_fd_sc_hd__decap_3 PHY_3148 ();
 sky130_fd_sc_hd__decap_3 PHY_3149 ();
 sky130_fd_sc_hd__decap_3 PHY_3150 ();
 sky130_fd_sc_hd__decap_3 PHY_3151 ();
 sky130_fd_sc_hd__decap_3 PHY_3152 ();
 sky130_fd_sc_hd__decap_3 PHY_3153 ();
 sky130_fd_sc_hd__decap_3 PHY_3154 ();
 sky130_fd_sc_hd__decap_3 PHY_3155 ();
 sky130_fd_sc_hd__decap_3 PHY_3156 ();
 sky130_fd_sc_hd__decap_3 PHY_3157 ();
 sky130_fd_sc_hd__decap_3 PHY_3158 ();
 sky130_fd_sc_hd__decap_3 PHY_3159 ();
 sky130_fd_sc_hd__decap_3 PHY_3160 ();
 sky130_fd_sc_hd__decap_3 PHY_3161 ();
 sky130_fd_sc_hd__decap_3 PHY_3162 ();
 sky130_fd_sc_hd__decap_3 PHY_3163 ();
 sky130_fd_sc_hd__decap_3 PHY_3164 ();
 sky130_fd_sc_hd__decap_3 PHY_3165 ();
 sky130_fd_sc_hd__decap_3 PHY_3166 ();
 sky130_fd_sc_hd__decap_3 PHY_3167 ();
 sky130_fd_sc_hd__decap_3 PHY_3168 ();
 sky130_fd_sc_hd__decap_3 PHY_3169 ();
 sky130_fd_sc_hd__decap_3 PHY_3170 ();
 sky130_fd_sc_hd__decap_3 PHY_3171 ();
 sky130_fd_sc_hd__decap_3 PHY_3172 ();
 sky130_fd_sc_hd__decap_3 PHY_3173 ();
 sky130_fd_sc_hd__decap_3 PHY_3174 ();
 sky130_fd_sc_hd__decap_3 PHY_3175 ();
 sky130_fd_sc_hd__decap_3 PHY_3176 ();
 sky130_fd_sc_hd__decap_3 PHY_3177 ();
 sky130_fd_sc_hd__decap_3 PHY_3178 ();
 sky130_fd_sc_hd__decap_3 PHY_3179 ();
 sky130_fd_sc_hd__decap_3 PHY_3180 ();
 sky130_fd_sc_hd__decap_3 PHY_3181 ();
 sky130_fd_sc_hd__decap_3 PHY_3182 ();
 sky130_fd_sc_hd__decap_3 PHY_3183 ();
 sky130_fd_sc_hd__decap_3 PHY_3184 ();
 sky130_fd_sc_hd__decap_3 PHY_3185 ();
 sky130_fd_sc_hd__decap_3 PHY_3186 ();
 sky130_fd_sc_hd__decap_3 PHY_3187 ();
 sky130_fd_sc_hd__decap_3 PHY_3188 ();
 sky130_fd_sc_hd__decap_3 PHY_3189 ();
 sky130_fd_sc_hd__decap_3 PHY_3190 ();
 sky130_fd_sc_hd__decap_3 PHY_3191 ();
 sky130_fd_sc_hd__decap_3 PHY_3192 ();
 sky130_fd_sc_hd__decap_3 PHY_3193 ();
 sky130_fd_sc_hd__decap_3 PHY_3194 ();
 sky130_fd_sc_hd__decap_3 PHY_3195 ();
 sky130_fd_sc_hd__decap_3 PHY_3196 ();
 sky130_fd_sc_hd__decap_3 PHY_3197 ();
 sky130_fd_sc_hd__decap_3 PHY_3198 ();
 sky130_fd_sc_hd__decap_3 PHY_3199 ();
 sky130_fd_sc_hd__decap_3 PHY_3200 ();
 sky130_fd_sc_hd__decap_3 PHY_3201 ();
 sky130_fd_sc_hd__decap_3 PHY_3202 ();
 sky130_fd_sc_hd__decap_3 PHY_3203 ();
 sky130_fd_sc_hd__decap_3 PHY_3204 ();
 sky130_fd_sc_hd__decap_3 PHY_3205 ();
 sky130_fd_sc_hd__decap_3 PHY_3206 ();
 sky130_fd_sc_hd__decap_3 PHY_3207 ();
 sky130_fd_sc_hd__decap_3 PHY_3208 ();
 sky130_fd_sc_hd__decap_3 PHY_3209 ();
 sky130_fd_sc_hd__decap_3 PHY_3210 ();
 sky130_fd_sc_hd__decap_3 PHY_3211 ();
 sky130_fd_sc_hd__decap_3 PHY_3212 ();
 sky130_fd_sc_hd__decap_3 PHY_3213 ();
 sky130_fd_sc_hd__decap_3 PHY_3214 ();
 sky130_fd_sc_hd__decap_3 PHY_3215 ();
 sky130_fd_sc_hd__decap_3 PHY_3216 ();
 sky130_fd_sc_hd__decap_3 PHY_3217 ();
 sky130_fd_sc_hd__decap_3 PHY_3218 ();
 sky130_fd_sc_hd__decap_3 PHY_3219 ();
 sky130_fd_sc_hd__decap_3 PHY_3220 ();
 sky130_fd_sc_hd__decap_3 PHY_3221 ();
 sky130_fd_sc_hd__decap_3 PHY_3222 ();
 sky130_fd_sc_hd__decap_3 PHY_3223 ();
 sky130_fd_sc_hd__decap_3 PHY_3224 ();
 sky130_fd_sc_hd__decap_3 PHY_3225 ();
 sky130_fd_sc_hd__decap_3 PHY_3226 ();
 sky130_fd_sc_hd__decap_3 PHY_3227 ();
 sky130_fd_sc_hd__decap_3 PHY_3228 ();
 sky130_fd_sc_hd__decap_3 PHY_3229 ();
 sky130_fd_sc_hd__decap_3 PHY_3230 ();
 sky130_fd_sc_hd__decap_3 PHY_3231 ();
 sky130_fd_sc_hd__decap_3 PHY_3232 ();
 sky130_fd_sc_hd__decap_3 PHY_3233 ();
 sky130_fd_sc_hd__decap_3 PHY_3234 ();
 sky130_fd_sc_hd__decap_3 PHY_3235 ();
 sky130_fd_sc_hd__decap_3 PHY_3236 ();
 sky130_fd_sc_hd__decap_3 PHY_3237 ();
 sky130_fd_sc_hd__decap_3 PHY_3238 ();
 sky130_fd_sc_hd__decap_3 PHY_3239 ();
 sky130_fd_sc_hd__decap_3 PHY_3240 ();
 sky130_fd_sc_hd__decap_3 PHY_3241 ();
 sky130_fd_sc_hd__decap_3 PHY_3242 ();
 sky130_fd_sc_hd__decap_3 PHY_3243 ();
 sky130_fd_sc_hd__decap_3 PHY_3244 ();
 sky130_fd_sc_hd__decap_3 PHY_3245 ();
 sky130_fd_sc_hd__decap_3 PHY_3246 ();
 sky130_fd_sc_hd__decap_3 PHY_3247 ();
 sky130_fd_sc_hd__decap_3 PHY_3248 ();
 sky130_fd_sc_hd__decap_3 PHY_3249 ();
 sky130_fd_sc_hd__decap_3 PHY_3250 ();
 sky130_fd_sc_hd__decap_3 PHY_3251 ();
 sky130_fd_sc_hd__decap_3 PHY_3252 ();
 sky130_fd_sc_hd__decap_3 PHY_3253 ();
 sky130_fd_sc_hd__decap_3 PHY_3254 ();
 sky130_fd_sc_hd__decap_3 PHY_3255 ();
 sky130_fd_sc_hd__decap_3 PHY_3256 ();
 sky130_fd_sc_hd__decap_3 PHY_3257 ();
 sky130_fd_sc_hd__decap_3 PHY_3258 ();
 sky130_fd_sc_hd__decap_3 PHY_3259 ();
 sky130_fd_sc_hd__decap_3 PHY_3260 ();
 sky130_fd_sc_hd__decap_3 PHY_3261 ();
 sky130_fd_sc_hd__decap_3 PHY_3262 ();
 sky130_fd_sc_hd__decap_3 PHY_3263 ();
 sky130_fd_sc_hd__decap_3 PHY_3264 ();
 sky130_fd_sc_hd__decap_3 PHY_3265 ();
 sky130_fd_sc_hd__decap_3 PHY_3266 ();
 sky130_fd_sc_hd__decap_3 PHY_3267 ();
 sky130_fd_sc_hd__decap_3 PHY_3268 ();
 sky130_fd_sc_hd__decap_3 PHY_3269 ();
 sky130_fd_sc_hd__decap_3 PHY_3270 ();
 sky130_fd_sc_hd__decap_3 PHY_3271 ();
 sky130_fd_sc_hd__decap_3 PHY_3272 ();
 sky130_fd_sc_hd__decap_3 PHY_3273 ();
 sky130_fd_sc_hd__decap_3 PHY_3274 ();
 sky130_fd_sc_hd__decap_3 PHY_3275 ();
 sky130_fd_sc_hd__decap_3 PHY_3276 ();
 sky130_fd_sc_hd__decap_3 PHY_3277 ();
 sky130_fd_sc_hd__decap_3 PHY_3278 ();
 sky130_fd_sc_hd__decap_3 PHY_3279 ();
 sky130_fd_sc_hd__decap_3 PHY_3280 ();
 sky130_fd_sc_hd__decap_3 PHY_3281 ();
 sky130_fd_sc_hd__decap_3 PHY_3282 ();
 sky130_fd_sc_hd__decap_3 PHY_3283 ();
 sky130_fd_sc_hd__decap_3 PHY_3284 ();
 sky130_fd_sc_hd__decap_3 PHY_3285 ();
 sky130_fd_sc_hd__decap_3 PHY_3286 ();
 sky130_fd_sc_hd__decap_3 PHY_3287 ();
 sky130_fd_sc_hd__decap_3 PHY_3288 ();
 sky130_fd_sc_hd__decap_3 PHY_3289 ();
 sky130_fd_sc_hd__decap_3 PHY_3290 ();
 sky130_fd_sc_hd__decap_3 PHY_3291 ();
 sky130_fd_sc_hd__decap_3 PHY_3292 ();
 sky130_fd_sc_hd__decap_3 PHY_3293 ();
 sky130_fd_sc_hd__decap_3 PHY_3294 ();
 sky130_fd_sc_hd__decap_3 PHY_3295 ();
 sky130_fd_sc_hd__decap_3 PHY_3296 ();
 sky130_fd_sc_hd__decap_3 PHY_3297 ();
 sky130_fd_sc_hd__decap_3 PHY_3298 ();
 sky130_fd_sc_hd__decap_3 PHY_3299 ();
 sky130_fd_sc_hd__decap_3 PHY_3300 ();
 sky130_fd_sc_hd__decap_3 PHY_3301 ();
 sky130_fd_sc_hd__decap_3 PHY_3302 ();
 sky130_fd_sc_hd__decap_3 PHY_3303 ();
 sky130_fd_sc_hd__decap_3 PHY_3304 ();
 sky130_fd_sc_hd__decap_3 PHY_3305 ();
 sky130_fd_sc_hd__decap_3 PHY_3306 ();
 sky130_fd_sc_hd__decap_3 PHY_3307 ();
 sky130_fd_sc_hd__decap_3 PHY_3308 ();
 sky130_fd_sc_hd__decap_3 PHY_3309 ();
 sky130_fd_sc_hd__decap_3 PHY_3310 ();
 sky130_fd_sc_hd__decap_3 PHY_3311 ();
 sky130_fd_sc_hd__decap_3 PHY_3312 ();
 sky130_fd_sc_hd__decap_3 PHY_3313 ();
 sky130_fd_sc_hd__decap_3 PHY_3314 ();
 sky130_fd_sc_hd__decap_3 PHY_3315 ();
 sky130_fd_sc_hd__decap_3 PHY_3316 ();
 sky130_fd_sc_hd__decap_3 PHY_3317 ();
 sky130_fd_sc_hd__decap_3 PHY_3318 ();
 sky130_fd_sc_hd__decap_3 PHY_3319 ();
 sky130_fd_sc_hd__decap_3 PHY_3320 ();
 sky130_fd_sc_hd__decap_3 PHY_3321 ();
 sky130_fd_sc_hd__decap_3 PHY_3322 ();
 sky130_fd_sc_hd__decap_3 PHY_3323 ();
 sky130_fd_sc_hd__decap_3 PHY_3324 ();
 sky130_fd_sc_hd__decap_3 PHY_3325 ();
 sky130_fd_sc_hd__decap_3 PHY_3326 ();
 sky130_fd_sc_hd__decap_3 PHY_3327 ();
 sky130_fd_sc_hd__decap_3 PHY_3328 ();
 sky130_fd_sc_hd__decap_3 PHY_3329 ();
 sky130_fd_sc_hd__decap_3 PHY_3330 ();
 sky130_fd_sc_hd__decap_3 PHY_3331 ();
 sky130_fd_sc_hd__decap_3 PHY_3332 ();
 sky130_fd_sc_hd__decap_3 PHY_3333 ();
 sky130_fd_sc_hd__decap_3 PHY_3334 ();
 sky130_fd_sc_hd__decap_3 PHY_3335 ();
 sky130_fd_sc_hd__decap_3 PHY_3336 ();
 sky130_fd_sc_hd__decap_3 PHY_3337 ();
 sky130_fd_sc_hd__decap_3 PHY_3338 ();
 sky130_fd_sc_hd__decap_3 PHY_3339 ();
 sky130_fd_sc_hd__decap_3 PHY_3340 ();
 sky130_fd_sc_hd__decap_3 PHY_3341 ();
 sky130_fd_sc_hd__decap_3 PHY_3342 ();
 sky130_fd_sc_hd__decap_3 PHY_3343 ();
 sky130_fd_sc_hd__decap_3 PHY_3344 ();
 sky130_fd_sc_hd__decap_3 PHY_3345 ();
 sky130_fd_sc_hd__decap_3 PHY_3346 ();
 sky130_fd_sc_hd__decap_3 PHY_3347 ();
 sky130_fd_sc_hd__decap_3 PHY_3348 ();
 sky130_fd_sc_hd__decap_3 PHY_3349 ();
 sky130_fd_sc_hd__decap_3 PHY_3350 ();
 sky130_fd_sc_hd__decap_3 PHY_3351 ();
 sky130_fd_sc_hd__decap_3 PHY_3352 ();
 sky130_fd_sc_hd__decap_3 PHY_3353 ();
 sky130_fd_sc_hd__decap_3 PHY_3354 ();
 sky130_fd_sc_hd__decap_3 PHY_3355 ();
 sky130_fd_sc_hd__decap_3 PHY_3356 ();
 sky130_fd_sc_hd__decap_3 PHY_3357 ();
 sky130_fd_sc_hd__decap_3 PHY_3358 ();
 sky130_fd_sc_hd__decap_3 PHY_3359 ();
 sky130_fd_sc_hd__decap_3 PHY_3360 ();
 sky130_fd_sc_hd__decap_3 PHY_3361 ();
 sky130_fd_sc_hd__decap_3 PHY_3362 ();
 sky130_fd_sc_hd__decap_3 PHY_3363 ();
 sky130_fd_sc_hd__decap_3 PHY_3364 ();
 sky130_fd_sc_hd__decap_3 PHY_3365 ();
 sky130_fd_sc_hd__decap_3 PHY_3366 ();
 sky130_fd_sc_hd__decap_3 PHY_3367 ();
 sky130_fd_sc_hd__decap_3 PHY_3368 ();
 sky130_fd_sc_hd__decap_3 PHY_3369 ();
 sky130_fd_sc_hd__decap_3 PHY_3370 ();
 sky130_fd_sc_hd__decap_3 PHY_3371 ();
 sky130_fd_sc_hd__decap_3 PHY_3372 ();
 sky130_fd_sc_hd__decap_3 PHY_3373 ();
 sky130_fd_sc_hd__decap_3 PHY_3374 ();
 sky130_fd_sc_hd__decap_3 PHY_3375 ();
 sky130_fd_sc_hd__decap_3 PHY_3376 ();
 sky130_fd_sc_hd__decap_3 PHY_3377 ();
 sky130_fd_sc_hd__decap_3 PHY_3378 ();
 sky130_fd_sc_hd__decap_3 PHY_3379 ();
 sky130_fd_sc_hd__decap_3 PHY_3380 ();
 sky130_fd_sc_hd__decap_3 PHY_3381 ();
 sky130_fd_sc_hd__decap_3 PHY_3382 ();
 sky130_fd_sc_hd__decap_3 PHY_3383 ();
 sky130_fd_sc_hd__decap_3 PHY_3384 ();
 sky130_fd_sc_hd__decap_3 PHY_3385 ();
 sky130_fd_sc_hd__decap_3 PHY_3386 ();
 sky130_fd_sc_hd__decap_3 PHY_3387 ();
 sky130_fd_sc_hd__decap_3 PHY_3388 ();
 sky130_fd_sc_hd__decap_3 PHY_3389 ();
 sky130_fd_sc_hd__decap_3 PHY_3390 ();
 sky130_fd_sc_hd__decap_3 PHY_3391 ();
 sky130_fd_sc_hd__decap_3 PHY_3392 ();
 sky130_fd_sc_hd__decap_3 PHY_3393 ();
 sky130_fd_sc_hd__decap_3 PHY_3394 ();
 sky130_fd_sc_hd__decap_3 PHY_3395 ();
 sky130_fd_sc_hd__decap_3 PHY_3396 ();
 sky130_fd_sc_hd__decap_3 PHY_3397 ();
 sky130_fd_sc_hd__decap_3 PHY_3398 ();
 sky130_fd_sc_hd__decap_3 PHY_3399 ();
 sky130_fd_sc_hd__decap_3 PHY_3400 ();
 sky130_fd_sc_hd__decap_3 PHY_3401 ();
 sky130_fd_sc_hd__decap_3 PHY_3402 ();
 sky130_fd_sc_hd__decap_3 PHY_3403 ();
 sky130_fd_sc_hd__decap_3 PHY_3404 ();
 sky130_fd_sc_hd__decap_3 PHY_3405 ();
 sky130_fd_sc_hd__decap_3 PHY_3406 ();
 sky130_fd_sc_hd__decap_3 PHY_3407 ();
 sky130_fd_sc_hd__decap_3 PHY_3408 ();
 sky130_fd_sc_hd__decap_3 PHY_3409 ();
 sky130_fd_sc_hd__decap_3 PHY_3410 ();
 sky130_fd_sc_hd__decap_3 PHY_3411 ();
 sky130_fd_sc_hd__decap_3 PHY_3412 ();
 sky130_fd_sc_hd__decap_3 PHY_3413 ();
 sky130_fd_sc_hd__decap_3 PHY_3414 ();
 sky130_fd_sc_hd__decap_3 PHY_3415 ();
 sky130_fd_sc_hd__decap_3 PHY_3416 ();
 sky130_fd_sc_hd__decap_3 PHY_3417 ();
 sky130_fd_sc_hd__decap_3 PHY_3418 ();
 sky130_fd_sc_hd__decap_3 PHY_3419 ();
 sky130_fd_sc_hd__decap_3 PHY_3420 ();
 sky130_fd_sc_hd__decap_3 PHY_3421 ();
 sky130_fd_sc_hd__decap_3 PHY_3422 ();
 sky130_fd_sc_hd__decap_3 PHY_3423 ();
 sky130_fd_sc_hd__decap_3 PHY_3424 ();
 sky130_fd_sc_hd__decap_3 PHY_3425 ();
 sky130_fd_sc_hd__decap_3 PHY_3426 ();
 sky130_fd_sc_hd__decap_3 PHY_3427 ();
 sky130_fd_sc_hd__decap_3 PHY_3428 ();
 sky130_fd_sc_hd__decap_3 PHY_3429 ();
 sky130_fd_sc_hd__decap_3 PHY_3430 ();
 sky130_fd_sc_hd__decap_3 PHY_3431 ();
 sky130_fd_sc_hd__decap_3 PHY_3432 ();
 sky130_fd_sc_hd__decap_3 PHY_3433 ();
 sky130_fd_sc_hd__decap_3 PHY_3434 ();
 sky130_fd_sc_hd__decap_3 PHY_3435 ();
 sky130_fd_sc_hd__decap_3 PHY_3436 ();
 sky130_fd_sc_hd__decap_3 PHY_3437 ();
 sky130_fd_sc_hd__decap_3 PHY_3438 ();
 sky130_fd_sc_hd__decap_3 PHY_3439 ();
 sky130_fd_sc_hd__decap_3 PHY_3440 ();
 sky130_fd_sc_hd__decap_3 PHY_3441 ();
 sky130_fd_sc_hd__decap_3 PHY_3442 ();
 sky130_fd_sc_hd__decap_3 PHY_3443 ();
 sky130_fd_sc_hd__decap_3 PHY_3444 ();
 sky130_fd_sc_hd__decap_3 PHY_3445 ();
 sky130_fd_sc_hd__decap_3 PHY_3446 ();
 sky130_fd_sc_hd__decap_3 PHY_3447 ();
 sky130_fd_sc_hd__decap_3 PHY_3448 ();
 sky130_fd_sc_hd__decap_3 PHY_3449 ();
 sky130_fd_sc_hd__decap_3 PHY_3450 ();
 sky130_fd_sc_hd__decap_3 PHY_3451 ();
 sky130_fd_sc_hd__decap_3 PHY_3452 ();
 sky130_fd_sc_hd__decap_3 PHY_3453 ();
 sky130_fd_sc_hd__decap_3 PHY_3454 ();
 sky130_fd_sc_hd__decap_3 PHY_3455 ();
 sky130_fd_sc_hd__decap_3 PHY_3456 ();
 sky130_fd_sc_hd__decap_3 PHY_3457 ();
 sky130_fd_sc_hd__decap_3 PHY_3458 ();
 sky130_fd_sc_hd__decap_3 PHY_3459 ();
 sky130_fd_sc_hd__decap_3 PHY_3460 ();
 sky130_fd_sc_hd__decap_3 PHY_3461 ();
 sky130_fd_sc_hd__decap_3 PHY_3462 ();
 sky130_fd_sc_hd__decap_3 PHY_3463 ();
 sky130_fd_sc_hd__decap_3 PHY_3464 ();
 sky130_fd_sc_hd__decap_3 PHY_3465 ();
 sky130_fd_sc_hd__decap_3 PHY_3466 ();
 sky130_fd_sc_hd__decap_3 PHY_3467 ();
 sky130_fd_sc_hd__decap_3 PHY_3468 ();
 sky130_fd_sc_hd__decap_3 PHY_3469 ();
 sky130_fd_sc_hd__decap_3 PHY_3470 ();
 sky130_fd_sc_hd__decap_3 PHY_3471 ();
 sky130_fd_sc_hd__decap_3 PHY_3472 ();
 sky130_fd_sc_hd__decap_3 PHY_3473 ();
 sky130_fd_sc_hd__decap_3 PHY_3474 ();
 sky130_fd_sc_hd__decap_3 PHY_3475 ();
 sky130_fd_sc_hd__decap_3 PHY_3476 ();
 sky130_fd_sc_hd__decap_3 PHY_3477 ();
 sky130_fd_sc_hd__decap_3 PHY_3478 ();
 sky130_fd_sc_hd__decap_3 PHY_3479 ();
 sky130_fd_sc_hd__decap_3 PHY_3480 ();
 sky130_fd_sc_hd__decap_3 PHY_3481 ();
 sky130_fd_sc_hd__decap_3 PHY_3482 ();
 sky130_fd_sc_hd__decap_3 PHY_3483 ();
 sky130_fd_sc_hd__decap_3 PHY_3484 ();
 sky130_fd_sc_hd__decap_3 PHY_3485 ();
 sky130_fd_sc_hd__decap_3 PHY_3486 ();
 sky130_fd_sc_hd__decap_3 PHY_3487 ();
 sky130_fd_sc_hd__decap_3 PHY_3488 ();
 sky130_fd_sc_hd__decap_3 PHY_3489 ();
 sky130_fd_sc_hd__decap_3 PHY_3490 ();
 sky130_fd_sc_hd__decap_3 PHY_3491 ();
 sky130_fd_sc_hd__decap_3 PHY_3492 ();
 sky130_fd_sc_hd__decap_3 PHY_3493 ();
 sky130_fd_sc_hd__decap_3 PHY_3494 ();
 sky130_fd_sc_hd__decap_3 PHY_3495 ();
 sky130_fd_sc_hd__decap_3 PHY_3496 ();
 sky130_fd_sc_hd__decap_3 PHY_3497 ();
 sky130_fd_sc_hd__decap_3 PHY_3498 ();
 sky130_fd_sc_hd__decap_3 PHY_3499 ();
 sky130_fd_sc_hd__decap_3 PHY_3500 ();
 sky130_fd_sc_hd__decap_3 PHY_3501 ();
 sky130_fd_sc_hd__decap_3 PHY_3502 ();
 sky130_fd_sc_hd__decap_3 PHY_3503 ();
 sky130_fd_sc_hd__decap_3 PHY_3504 ();
 sky130_fd_sc_hd__decap_3 PHY_3505 ();
 sky130_fd_sc_hd__decap_3 PHY_3506 ();
 sky130_fd_sc_hd__decap_3 PHY_3507 ();
 sky130_fd_sc_hd__decap_3 PHY_3508 ();
 sky130_fd_sc_hd__decap_3 PHY_3509 ();
 sky130_fd_sc_hd__decap_3 PHY_3510 ();
 sky130_fd_sc_hd__decap_3 PHY_3511 ();
 sky130_fd_sc_hd__decap_3 PHY_3512 ();
 sky130_fd_sc_hd__decap_3 PHY_3513 ();
 sky130_fd_sc_hd__decap_3 PHY_3514 ();
 sky130_fd_sc_hd__decap_3 PHY_3515 ();
 sky130_fd_sc_hd__decap_3 PHY_3516 ();
 sky130_fd_sc_hd__decap_3 PHY_3517 ();
 sky130_fd_sc_hd__decap_3 PHY_3518 ();
 sky130_fd_sc_hd__decap_3 PHY_3519 ();
 sky130_fd_sc_hd__decap_3 PHY_3520 ();
 sky130_fd_sc_hd__decap_3 PHY_3521 ();
 sky130_fd_sc_hd__decap_3 PHY_3522 ();
 sky130_fd_sc_hd__decap_3 PHY_3523 ();
 sky130_fd_sc_hd__decap_3 PHY_3524 ();
 sky130_fd_sc_hd__decap_3 PHY_3525 ();
 sky130_fd_sc_hd__decap_3 PHY_3526 ();
 sky130_fd_sc_hd__decap_3 PHY_3527 ();
 sky130_fd_sc_hd__decap_3 PHY_3528 ();
 sky130_fd_sc_hd__decap_3 PHY_3529 ();
 sky130_fd_sc_hd__decap_3 PHY_3530 ();
 sky130_fd_sc_hd__decap_3 PHY_3531 ();
 sky130_fd_sc_hd__decap_3 PHY_3532 ();
 sky130_fd_sc_hd__decap_3 PHY_3533 ();
 sky130_fd_sc_hd__decap_3 PHY_3534 ();
 sky130_fd_sc_hd__decap_3 PHY_3535 ();
 sky130_fd_sc_hd__decap_3 PHY_3536 ();
 sky130_fd_sc_hd__decap_3 PHY_3537 ();
 sky130_fd_sc_hd__decap_3 PHY_3538 ();
 sky130_fd_sc_hd__decap_3 PHY_3539 ();
 sky130_fd_sc_hd__decap_3 PHY_3540 ();
 sky130_fd_sc_hd__decap_3 PHY_3541 ();
 sky130_fd_sc_hd__decap_3 PHY_3542 ();
 sky130_fd_sc_hd__decap_3 PHY_3543 ();
 sky130_fd_sc_hd__decap_3 PHY_3544 ();
 sky130_fd_sc_hd__decap_3 PHY_3545 ();
 sky130_fd_sc_hd__decap_3 PHY_3546 ();
 sky130_fd_sc_hd__decap_3 PHY_3547 ();
 sky130_fd_sc_hd__decap_3 PHY_3548 ();
 sky130_fd_sc_hd__decap_3 PHY_3549 ();
 sky130_fd_sc_hd__decap_3 PHY_3550 ();
 sky130_fd_sc_hd__decap_3 PHY_3551 ();
 sky130_fd_sc_hd__decap_3 PHY_3552 ();
 sky130_fd_sc_hd__decap_3 PHY_3553 ();
 sky130_fd_sc_hd__decap_3 PHY_3554 ();
 sky130_fd_sc_hd__decap_3 PHY_3555 ();
 sky130_fd_sc_hd__decap_3 PHY_3556 ();
 sky130_fd_sc_hd__decap_3 PHY_3557 ();
 sky130_fd_sc_hd__decap_3 PHY_3558 ();
 sky130_fd_sc_hd__decap_3 PHY_3559 ();
 sky130_fd_sc_hd__decap_3 PHY_3560 ();
 sky130_fd_sc_hd__decap_3 PHY_3561 ();
 sky130_fd_sc_hd__decap_3 PHY_3562 ();
 sky130_fd_sc_hd__decap_3 PHY_3563 ();
 sky130_fd_sc_hd__decap_3 PHY_3564 ();
 sky130_fd_sc_hd__decap_3 PHY_3565 ();
 sky130_fd_sc_hd__decap_3 PHY_3566 ();
 sky130_fd_sc_hd__decap_3 PHY_3567 ();
 sky130_fd_sc_hd__decap_3 PHY_3568 ();
 sky130_fd_sc_hd__decap_3 PHY_3569 ();
 sky130_fd_sc_hd__decap_3 PHY_3570 ();
 sky130_fd_sc_hd__decap_3 PHY_3571 ();
 sky130_fd_sc_hd__decap_3 PHY_3572 ();
 sky130_fd_sc_hd__decap_3 PHY_3573 ();
 sky130_fd_sc_hd__decap_3 PHY_3574 ();
 sky130_fd_sc_hd__decap_3 PHY_3575 ();
 sky130_fd_sc_hd__decap_3 PHY_3576 ();
 sky130_fd_sc_hd__decap_3 PHY_3577 ();
 sky130_fd_sc_hd__decap_3 PHY_3578 ();
 sky130_fd_sc_hd__decap_3 PHY_3579 ();
 sky130_fd_sc_hd__decap_3 PHY_3580 ();
 sky130_fd_sc_hd__decap_3 PHY_3581 ();
 sky130_fd_sc_hd__decap_3 PHY_3582 ();
 sky130_fd_sc_hd__decap_3 PHY_3583 ();
 sky130_fd_sc_hd__decap_3 PHY_3584 ();
 sky130_fd_sc_hd__decap_3 PHY_3585 ();
 sky130_fd_sc_hd__decap_3 PHY_3586 ();
 sky130_fd_sc_hd__decap_3 PHY_3587 ();
 sky130_fd_sc_hd__decap_3 PHY_3588 ();
 sky130_fd_sc_hd__decap_3 PHY_3589 ();
 sky130_fd_sc_hd__decap_3 PHY_3590 ();
 sky130_fd_sc_hd__decap_3 PHY_3591 ();
 sky130_fd_sc_hd__decap_3 PHY_3592 ();
 sky130_fd_sc_hd__decap_3 PHY_3593 ();
 sky130_fd_sc_hd__decap_3 PHY_3594 ();
 sky130_fd_sc_hd__decap_3 PHY_3595 ();
 sky130_fd_sc_hd__decap_3 PHY_3596 ();
 sky130_fd_sc_hd__decap_3 PHY_3597 ();
 sky130_fd_sc_hd__decap_3 PHY_3598 ();
 sky130_fd_sc_hd__decap_3 PHY_3599 ();
 sky130_fd_sc_hd__decap_3 PHY_3600 ();
 sky130_fd_sc_hd__decap_3 PHY_3601 ();
 sky130_fd_sc_hd__decap_3 PHY_3602 ();
 sky130_fd_sc_hd__decap_3 PHY_3603 ();
 sky130_fd_sc_hd__decap_3 PHY_3604 ();
 sky130_fd_sc_hd__decap_3 PHY_3605 ();
 sky130_fd_sc_hd__decap_3 PHY_3606 ();
 sky130_fd_sc_hd__decap_3 PHY_3607 ();
 sky130_fd_sc_hd__decap_3 PHY_3608 ();
 sky130_fd_sc_hd__decap_3 PHY_3609 ();
 sky130_fd_sc_hd__decap_3 PHY_3610 ();
 sky130_fd_sc_hd__decap_3 PHY_3611 ();
 sky130_fd_sc_hd__decap_3 PHY_3612 ();
 sky130_fd_sc_hd__decap_3 PHY_3613 ();
 sky130_fd_sc_hd__decap_3 PHY_3614 ();
 sky130_fd_sc_hd__decap_3 PHY_3615 ();
 sky130_fd_sc_hd__decap_3 PHY_3616 ();
 sky130_fd_sc_hd__decap_3 PHY_3617 ();
 sky130_fd_sc_hd__decap_3 PHY_3618 ();
 sky130_fd_sc_hd__decap_3 PHY_3619 ();
 sky130_fd_sc_hd__decap_3 PHY_3620 ();
 sky130_fd_sc_hd__decap_3 PHY_3621 ();
 sky130_fd_sc_hd__decap_3 PHY_3622 ();
 sky130_fd_sc_hd__decap_3 PHY_3623 ();
 sky130_fd_sc_hd__decap_3 PHY_3624 ();
 sky130_fd_sc_hd__decap_3 PHY_3625 ();
 sky130_fd_sc_hd__decap_3 PHY_3626 ();
 sky130_fd_sc_hd__decap_3 PHY_3627 ();
 sky130_fd_sc_hd__decap_3 PHY_3628 ();
 sky130_fd_sc_hd__decap_3 PHY_3629 ();
 sky130_fd_sc_hd__decap_3 PHY_3630 ();
 sky130_fd_sc_hd__decap_3 PHY_3631 ();
 sky130_fd_sc_hd__decap_3 PHY_3632 ();
 sky130_fd_sc_hd__decap_3 PHY_3633 ();
 sky130_fd_sc_hd__decap_3 PHY_3634 ();
 sky130_fd_sc_hd__decap_3 PHY_3635 ();
 sky130_fd_sc_hd__decap_3 PHY_3636 ();
 sky130_fd_sc_hd__decap_3 PHY_3637 ();
 sky130_fd_sc_hd__decap_3 PHY_3638 ();
 sky130_fd_sc_hd__decap_3 PHY_3639 ();
 sky130_fd_sc_hd__decap_3 PHY_3640 ();
 sky130_fd_sc_hd__decap_3 PHY_3641 ();
 sky130_fd_sc_hd__decap_3 PHY_3642 ();
 sky130_fd_sc_hd__decap_3 PHY_3643 ();
 sky130_fd_sc_hd__decap_3 PHY_3644 ();
 sky130_fd_sc_hd__decap_3 PHY_3645 ();
 sky130_fd_sc_hd__decap_3 PHY_3646 ();
 sky130_fd_sc_hd__decap_3 PHY_3647 ();
 sky130_fd_sc_hd__decap_3 PHY_3648 ();
 sky130_fd_sc_hd__decap_3 PHY_3649 ();
 sky130_fd_sc_hd__decap_3 PHY_3650 ();
 sky130_fd_sc_hd__decap_3 PHY_3651 ();
 sky130_fd_sc_hd__decap_3 PHY_3652 ();
 sky130_fd_sc_hd__decap_3 PHY_3653 ();
 sky130_fd_sc_hd__decap_3 PHY_3654 ();
 sky130_fd_sc_hd__decap_3 PHY_3655 ();
 sky130_fd_sc_hd__decap_3 PHY_3656 ();
 sky130_fd_sc_hd__decap_3 PHY_3657 ();
 sky130_fd_sc_hd__decap_3 PHY_3658 ();
 sky130_fd_sc_hd__decap_3 PHY_3659 ();
 sky130_fd_sc_hd__decap_3 PHY_3660 ();
 sky130_fd_sc_hd__decap_3 PHY_3661 ();
 sky130_fd_sc_hd__decap_3 PHY_3662 ();
 sky130_fd_sc_hd__decap_3 PHY_3663 ();
 sky130_fd_sc_hd__decap_3 PHY_3664 ();
 sky130_fd_sc_hd__decap_3 PHY_3665 ();
 sky130_fd_sc_hd__decap_3 PHY_3666 ();
 sky130_fd_sc_hd__decap_3 PHY_3667 ();
 sky130_fd_sc_hd__decap_3 PHY_3668 ();
 sky130_fd_sc_hd__decap_3 PHY_3669 ();
 sky130_fd_sc_hd__decap_3 PHY_3670 ();
 sky130_fd_sc_hd__decap_3 PHY_3671 ();
 sky130_fd_sc_hd__decap_3 PHY_3672 ();
 sky130_fd_sc_hd__decap_3 PHY_3673 ();
 sky130_fd_sc_hd__decap_3 PHY_3674 ();
 sky130_fd_sc_hd__decap_3 PHY_3675 ();
 sky130_fd_sc_hd__decap_3 PHY_3676 ();
 sky130_fd_sc_hd__decap_3 PHY_3677 ();
 sky130_fd_sc_hd__decap_3 PHY_3678 ();
 sky130_fd_sc_hd__decap_3 PHY_3679 ();
 sky130_fd_sc_hd__decap_3 PHY_3680 ();
 sky130_fd_sc_hd__decap_3 PHY_3681 ();
 sky130_fd_sc_hd__decap_3 PHY_3682 ();
 sky130_fd_sc_hd__decap_3 PHY_3683 ();
 sky130_fd_sc_hd__decap_3 PHY_3684 ();
 sky130_fd_sc_hd__decap_3 PHY_3685 ();
 sky130_fd_sc_hd__decap_3 PHY_3686 ();
 sky130_fd_sc_hd__decap_3 PHY_3687 ();
 sky130_fd_sc_hd__decap_3 PHY_3688 ();
 sky130_fd_sc_hd__decap_3 PHY_3689 ();
 sky130_fd_sc_hd__decap_3 PHY_3690 ();
 sky130_fd_sc_hd__decap_3 PHY_3691 ();
 sky130_fd_sc_hd__decap_3 PHY_3692 ();
 sky130_fd_sc_hd__decap_3 PHY_3693 ();
 sky130_fd_sc_hd__decap_3 PHY_3694 ();
 sky130_fd_sc_hd__decap_3 PHY_3695 ();
 sky130_fd_sc_hd__decap_3 PHY_3696 ();
 sky130_fd_sc_hd__decap_3 PHY_3697 ();
 sky130_fd_sc_hd__decap_3 PHY_3698 ();
 sky130_fd_sc_hd__decap_3 PHY_3699 ();
 sky130_fd_sc_hd__decap_3 PHY_3700 ();
 sky130_fd_sc_hd__decap_3 PHY_3701 ();
 sky130_fd_sc_hd__decap_3 PHY_3702 ();
 sky130_fd_sc_hd__decap_3 PHY_3703 ();
 sky130_fd_sc_hd__decap_3 PHY_3704 ();
 sky130_fd_sc_hd__decap_3 PHY_3705 ();
 sky130_fd_sc_hd__decap_3 PHY_3706 ();
 sky130_fd_sc_hd__decap_3 PHY_3707 ();
 sky130_fd_sc_hd__decap_3 PHY_3708 ();
 sky130_fd_sc_hd__decap_3 PHY_3709 ();
 sky130_fd_sc_hd__decap_3 PHY_3710 ();
 sky130_fd_sc_hd__decap_3 PHY_3711 ();
 sky130_fd_sc_hd__decap_3 PHY_3712 ();
 sky130_fd_sc_hd__decap_3 PHY_3713 ();
 sky130_fd_sc_hd__decap_3 PHY_3714 ();
 sky130_fd_sc_hd__decap_3 PHY_3715 ();
 sky130_fd_sc_hd__decap_3 PHY_3716 ();
 sky130_fd_sc_hd__decap_3 PHY_3717 ();
 sky130_fd_sc_hd__decap_3 PHY_3718 ();
 sky130_fd_sc_hd__decap_3 PHY_3719 ();
 sky130_fd_sc_hd__decap_3 PHY_3720 ();
 sky130_fd_sc_hd__decap_3 PHY_3721 ();
 sky130_fd_sc_hd__decap_3 PHY_3722 ();
 sky130_fd_sc_hd__decap_3 PHY_3723 ();
 sky130_fd_sc_hd__decap_3 PHY_3724 ();
 sky130_fd_sc_hd__decap_3 PHY_3725 ();
 sky130_fd_sc_hd__decap_3 PHY_3726 ();
 sky130_fd_sc_hd__decap_3 PHY_3727 ();
 sky130_fd_sc_hd__decap_3 PHY_3728 ();
 sky130_fd_sc_hd__decap_3 PHY_3729 ();
 sky130_fd_sc_hd__decap_3 PHY_3730 ();
 sky130_fd_sc_hd__decap_3 PHY_3731 ();
 sky130_fd_sc_hd__decap_3 PHY_3732 ();
 sky130_fd_sc_hd__decap_3 PHY_3733 ();
 sky130_fd_sc_hd__decap_3 PHY_3734 ();
 sky130_fd_sc_hd__decap_3 PHY_3735 ();
 sky130_fd_sc_hd__decap_3 PHY_3736 ();
 sky130_fd_sc_hd__decap_3 PHY_3737 ();
 sky130_fd_sc_hd__decap_3 PHY_3738 ();
 sky130_fd_sc_hd__decap_3 PHY_3739 ();
 sky130_fd_sc_hd__decap_3 PHY_3740 ();
 sky130_fd_sc_hd__decap_3 PHY_3741 ();
 sky130_fd_sc_hd__decap_3 PHY_3742 ();
 sky130_fd_sc_hd__decap_3 PHY_3743 ();
 sky130_fd_sc_hd__decap_3 PHY_3744 ();
 sky130_fd_sc_hd__decap_3 PHY_3745 ();
 sky130_fd_sc_hd__decap_3 PHY_3746 ();
 sky130_fd_sc_hd__decap_3 PHY_3747 ();
 sky130_fd_sc_hd__decap_3 PHY_3748 ();
 sky130_fd_sc_hd__decap_3 PHY_3749 ();
 sky130_fd_sc_hd__decap_3 PHY_3750 ();
 sky130_fd_sc_hd__decap_3 PHY_3751 ();
 sky130_fd_sc_hd__decap_3 PHY_3752 ();
 sky130_fd_sc_hd__decap_3 PHY_3753 ();
 sky130_fd_sc_hd__decap_3 PHY_3754 ();
 sky130_fd_sc_hd__decap_3 PHY_3755 ();
 sky130_fd_sc_hd__decap_3 PHY_3756 ();
 sky130_fd_sc_hd__decap_3 PHY_3757 ();
 sky130_fd_sc_hd__decap_3 PHY_3758 ();
 sky130_fd_sc_hd__decap_3 PHY_3759 ();
 sky130_fd_sc_hd__decap_3 PHY_3760 ();
 sky130_fd_sc_hd__decap_3 PHY_3761 ();
 sky130_fd_sc_hd__decap_3 PHY_3762 ();
 sky130_fd_sc_hd__decap_3 PHY_3763 ();
 sky130_fd_sc_hd__decap_3 PHY_3764 ();
 sky130_fd_sc_hd__decap_3 PHY_3765 ();
 sky130_fd_sc_hd__decap_3 PHY_3766 ();
 sky130_fd_sc_hd__decap_3 PHY_3767 ();
 sky130_fd_sc_hd__decap_3 PHY_3768 ();
 sky130_fd_sc_hd__decap_3 PHY_3769 ();
 sky130_fd_sc_hd__decap_3 PHY_3770 ();
 sky130_fd_sc_hd__decap_3 PHY_3771 ();
 sky130_fd_sc_hd__decap_3 PHY_3772 ();
 sky130_fd_sc_hd__decap_3 PHY_3773 ();
 sky130_fd_sc_hd__decap_3 PHY_3774 ();
 sky130_fd_sc_hd__decap_3 PHY_3775 ();
 sky130_fd_sc_hd__decap_3 PHY_3776 ();
 sky130_fd_sc_hd__decap_3 PHY_3777 ();
 sky130_fd_sc_hd__decap_3 PHY_3778 ();
 sky130_fd_sc_hd__decap_3 PHY_3779 ();
 sky130_fd_sc_hd__decap_3 PHY_3780 ();
 sky130_fd_sc_hd__decap_3 PHY_3781 ();
 sky130_fd_sc_hd__decap_3 PHY_3782 ();
 sky130_fd_sc_hd__decap_3 PHY_3783 ();
 sky130_fd_sc_hd__decap_3 PHY_3784 ();
 sky130_fd_sc_hd__decap_3 PHY_3785 ();
 sky130_fd_sc_hd__decap_3 PHY_3786 ();
 sky130_fd_sc_hd__decap_3 PHY_3787 ();
 sky130_fd_sc_hd__decap_3 PHY_3788 ();
 sky130_fd_sc_hd__decap_3 PHY_3789 ();
 sky130_fd_sc_hd__decap_3 PHY_3790 ();
 sky130_fd_sc_hd__decap_3 PHY_3791 ();
 sky130_fd_sc_hd__decap_3 PHY_3792 ();
 sky130_fd_sc_hd__decap_3 PHY_3793 ();
 sky130_fd_sc_hd__decap_3 PHY_3794 ();
 sky130_fd_sc_hd__decap_3 PHY_3795 ();
 sky130_fd_sc_hd__decap_3 PHY_3796 ();
 sky130_fd_sc_hd__decap_3 PHY_3797 ();
 sky130_fd_sc_hd__decap_3 PHY_3798 ();
 sky130_fd_sc_hd__decap_3 PHY_3799 ();
 sky130_fd_sc_hd__decap_3 PHY_3800 ();
 sky130_fd_sc_hd__decap_3 PHY_3801 ();
 sky130_fd_sc_hd__decap_3 PHY_3802 ();
 sky130_fd_sc_hd__decap_3 PHY_3803 ();
 sky130_fd_sc_hd__decap_3 PHY_3804 ();
 sky130_fd_sc_hd__decap_3 PHY_3805 ();
 sky130_fd_sc_hd__decap_3 PHY_3806 ();
 sky130_fd_sc_hd__decap_3 PHY_3807 ();
 sky130_fd_sc_hd__decap_3 PHY_3808 ();
 sky130_fd_sc_hd__decap_3 PHY_3809 ();
 sky130_fd_sc_hd__decap_3 PHY_3810 ();
 sky130_fd_sc_hd__decap_3 PHY_3811 ();
 sky130_fd_sc_hd__decap_3 PHY_3812 ();
 sky130_fd_sc_hd__decap_3 PHY_3813 ();
 sky130_fd_sc_hd__decap_3 PHY_3814 ();
 sky130_fd_sc_hd__decap_3 PHY_3815 ();
 sky130_fd_sc_hd__decap_3 PHY_3816 ();
 sky130_fd_sc_hd__decap_3 PHY_3817 ();
 sky130_fd_sc_hd__decap_3 PHY_3818 ();
 sky130_fd_sc_hd__decap_3 PHY_3819 ();
 sky130_fd_sc_hd__decap_3 PHY_3820 ();
 sky130_fd_sc_hd__decap_3 PHY_3821 ();
 sky130_fd_sc_hd__decap_3 PHY_3822 ();
 sky130_fd_sc_hd__decap_3 PHY_3823 ();
 sky130_fd_sc_hd__decap_3 PHY_3824 ();
 sky130_fd_sc_hd__decap_3 PHY_3825 ();
 sky130_fd_sc_hd__decap_3 PHY_3826 ();
 sky130_fd_sc_hd__decap_3 PHY_3827 ();
 sky130_fd_sc_hd__decap_3 PHY_3828 ();
 sky130_fd_sc_hd__decap_3 PHY_3829 ();
 sky130_fd_sc_hd__decap_3 PHY_3830 ();
 sky130_fd_sc_hd__decap_3 PHY_3831 ();
 sky130_fd_sc_hd__decap_3 PHY_3832 ();
 sky130_fd_sc_hd__decap_3 PHY_3833 ();
 sky130_fd_sc_hd__decap_3 PHY_3834 ();
 sky130_fd_sc_hd__decap_3 PHY_3835 ();
 sky130_fd_sc_hd__decap_3 PHY_3836 ();
 sky130_fd_sc_hd__decap_3 PHY_3837 ();
 sky130_fd_sc_hd__decap_3 PHY_3838 ();
 sky130_fd_sc_hd__decap_3 PHY_3839 ();
 sky130_fd_sc_hd__decap_3 PHY_3840 ();
 sky130_fd_sc_hd__decap_3 PHY_3841 ();
 sky130_fd_sc_hd__decap_3 PHY_3842 ();
 sky130_fd_sc_hd__decap_3 PHY_3843 ();
 sky130_fd_sc_hd__decap_3 PHY_3844 ();
 sky130_fd_sc_hd__decap_3 PHY_3845 ();
 sky130_fd_sc_hd__decap_3 PHY_3846 ();
 sky130_fd_sc_hd__decap_3 PHY_3847 ();
 sky130_fd_sc_hd__decap_3 PHY_3848 ();
 sky130_fd_sc_hd__decap_3 PHY_3849 ();
 sky130_fd_sc_hd__decap_3 PHY_3850 ();
 sky130_fd_sc_hd__decap_3 PHY_3851 ();
 sky130_fd_sc_hd__decap_3 PHY_3852 ();
 sky130_fd_sc_hd__decap_3 PHY_3853 ();
 sky130_fd_sc_hd__decap_3 PHY_3854 ();
 sky130_fd_sc_hd__decap_3 PHY_3855 ();
 sky130_fd_sc_hd__decap_3 PHY_3856 ();
 sky130_fd_sc_hd__decap_3 PHY_3857 ();
 sky130_fd_sc_hd__decap_3 PHY_3858 ();
 sky130_fd_sc_hd__decap_3 PHY_3859 ();
 sky130_fd_sc_hd__decap_3 PHY_3860 ();
 sky130_fd_sc_hd__decap_3 PHY_3861 ();
 sky130_fd_sc_hd__decap_3 PHY_3862 ();
 sky130_fd_sc_hd__decap_3 PHY_3863 ();
 sky130_fd_sc_hd__decap_3 PHY_3864 ();
 sky130_fd_sc_hd__decap_3 PHY_3865 ();
 sky130_fd_sc_hd__decap_3 PHY_3866 ();
 sky130_fd_sc_hd__decap_3 PHY_3867 ();
 sky130_fd_sc_hd__decap_3 PHY_3868 ();
 sky130_fd_sc_hd__decap_3 PHY_3869 ();
 sky130_fd_sc_hd__decap_3 PHY_3870 ();
 sky130_fd_sc_hd__decap_3 PHY_3871 ();
 sky130_fd_sc_hd__decap_3 PHY_3872 ();
 sky130_fd_sc_hd__decap_3 PHY_3873 ();
 sky130_fd_sc_hd__decap_3 PHY_3874 ();
 sky130_fd_sc_hd__decap_3 PHY_3875 ();
 sky130_fd_sc_hd__decap_3 PHY_3876 ();
 sky130_fd_sc_hd__decap_3 PHY_3877 ();
 sky130_fd_sc_hd__decap_3 PHY_3878 ();
 sky130_fd_sc_hd__decap_3 PHY_3879 ();
 sky130_fd_sc_hd__decap_3 PHY_3880 ();
 sky130_fd_sc_hd__decap_3 PHY_3881 ();
 sky130_fd_sc_hd__decap_3 PHY_3882 ();
 sky130_fd_sc_hd__decap_3 PHY_3883 ();
 sky130_fd_sc_hd__decap_3 PHY_3884 ();
 sky130_fd_sc_hd__decap_3 PHY_3885 ();
 sky130_fd_sc_hd__decap_3 PHY_3886 ();
 sky130_fd_sc_hd__decap_3 PHY_3887 ();
 sky130_fd_sc_hd__decap_3 PHY_3888 ();
 sky130_fd_sc_hd__decap_3 PHY_3889 ();
 sky130_fd_sc_hd__decap_3 PHY_3890 ();
 sky130_fd_sc_hd__decap_3 PHY_3891 ();
 sky130_fd_sc_hd__decap_3 PHY_3892 ();
 sky130_fd_sc_hd__decap_3 PHY_3893 ();
 sky130_fd_sc_hd__decap_3 PHY_3894 ();
 sky130_fd_sc_hd__decap_3 PHY_3895 ();
 sky130_fd_sc_hd__decap_3 PHY_3896 ();
 sky130_fd_sc_hd__decap_3 PHY_3897 ();
 sky130_fd_sc_hd__decap_3 PHY_3898 ();
 sky130_fd_sc_hd__decap_3 PHY_3899 ();
 sky130_fd_sc_hd__decap_3 PHY_3900 ();
 sky130_fd_sc_hd__decap_3 PHY_3901 ();
 sky130_fd_sc_hd__decap_3 PHY_3902 ();
 sky130_fd_sc_hd__decap_3 PHY_3903 ();
 sky130_fd_sc_hd__decap_3 PHY_3904 ();
 sky130_fd_sc_hd__decap_3 PHY_3905 ();
 sky130_fd_sc_hd__decap_3 PHY_3906 ();
 sky130_fd_sc_hd__decap_3 PHY_3907 ();
 sky130_fd_sc_hd__decap_3 PHY_3908 ();
 sky130_fd_sc_hd__decap_3 PHY_3909 ();
 sky130_fd_sc_hd__decap_3 PHY_3910 ();
 sky130_fd_sc_hd__decap_3 PHY_3911 ();
 sky130_fd_sc_hd__decap_3 PHY_3912 ();
 sky130_fd_sc_hd__decap_3 PHY_3913 ();
 sky130_fd_sc_hd__decap_3 PHY_3914 ();
 sky130_fd_sc_hd__decap_3 PHY_3915 ();
 sky130_fd_sc_hd__decap_3 PHY_3916 ();
 sky130_fd_sc_hd__decap_3 PHY_3917 ();
 sky130_fd_sc_hd__decap_3 PHY_3918 ();
 sky130_fd_sc_hd__decap_3 PHY_3919 ();
 sky130_fd_sc_hd__decap_3 PHY_3920 ();
 sky130_fd_sc_hd__decap_3 PHY_3921 ();
 sky130_fd_sc_hd__decap_3 PHY_3922 ();
 sky130_fd_sc_hd__decap_3 PHY_3923 ();
 sky130_fd_sc_hd__decap_3 PHY_3924 ();
 sky130_fd_sc_hd__decap_3 PHY_3925 ();
 sky130_fd_sc_hd__decap_3 PHY_3926 ();
 sky130_fd_sc_hd__decap_3 PHY_3927 ();
 sky130_fd_sc_hd__decap_3 PHY_3928 ();
 sky130_fd_sc_hd__decap_3 PHY_3929 ();
 sky130_fd_sc_hd__decap_3 PHY_3930 ();
 sky130_fd_sc_hd__decap_3 PHY_3931 ();
 sky130_fd_sc_hd__decap_3 PHY_3932 ();
 sky130_fd_sc_hd__decap_3 PHY_3933 ();
 sky130_fd_sc_hd__decap_3 PHY_3934 ();
 sky130_fd_sc_hd__decap_3 PHY_3935 ();
 sky130_fd_sc_hd__decap_3 PHY_3936 ();
 sky130_fd_sc_hd__decap_3 PHY_3937 ();
 sky130_fd_sc_hd__decap_3 PHY_3938 ();
 sky130_fd_sc_hd__decap_3 PHY_3939 ();
 sky130_fd_sc_hd__decap_3 PHY_3940 ();
 sky130_fd_sc_hd__decap_3 PHY_3941 ();
 sky130_fd_sc_hd__decap_3 PHY_3942 ();
 sky130_fd_sc_hd__decap_3 PHY_3943 ();
 sky130_fd_sc_hd__decap_3 PHY_3944 ();
 sky130_fd_sc_hd__decap_3 PHY_3945 ();
 sky130_fd_sc_hd__decap_3 PHY_3946 ();
 sky130_fd_sc_hd__decap_3 PHY_3947 ();
 sky130_fd_sc_hd__decap_3 PHY_3948 ();
 sky130_fd_sc_hd__decap_3 PHY_3949 ();
 sky130_fd_sc_hd__decap_3 PHY_3950 ();
 sky130_fd_sc_hd__decap_3 PHY_3951 ();
 sky130_fd_sc_hd__decap_3 PHY_3952 ();
 sky130_fd_sc_hd__decap_3 PHY_3953 ();
 sky130_fd_sc_hd__decap_3 PHY_3954 ();
 sky130_fd_sc_hd__decap_3 PHY_3955 ();
 sky130_fd_sc_hd__decap_3 PHY_3956 ();
 sky130_fd_sc_hd__decap_3 PHY_3957 ();
 sky130_fd_sc_hd__decap_3 PHY_3958 ();
 sky130_fd_sc_hd__decap_3 PHY_3959 ();
 sky130_fd_sc_hd__decap_3 PHY_3960 ();
 sky130_fd_sc_hd__decap_3 PHY_3961 ();
 sky130_fd_sc_hd__decap_3 PHY_3962 ();
 sky130_fd_sc_hd__decap_3 PHY_3963 ();
 sky130_fd_sc_hd__decap_3 PHY_3964 ();
 sky130_fd_sc_hd__decap_3 PHY_3965 ();
 sky130_fd_sc_hd__decap_3 PHY_3966 ();
 sky130_fd_sc_hd__decap_3 PHY_3967 ();
 sky130_fd_sc_hd__decap_3 PHY_3968 ();
 sky130_fd_sc_hd__decap_3 PHY_3969 ();
 sky130_fd_sc_hd__decap_3 PHY_3970 ();
 sky130_fd_sc_hd__decap_3 PHY_3971 ();
 sky130_fd_sc_hd__decap_3 PHY_3972 ();
 sky130_fd_sc_hd__decap_3 PHY_3973 ();
 sky130_fd_sc_hd__decap_3 PHY_3974 ();
 sky130_fd_sc_hd__decap_3 PHY_3975 ();
 sky130_fd_sc_hd__decap_3 PHY_3976 ();
 sky130_fd_sc_hd__decap_3 PHY_3977 ();
 sky130_fd_sc_hd__decap_3 PHY_3978 ();
 sky130_fd_sc_hd__decap_3 PHY_3979 ();
 sky130_fd_sc_hd__decap_3 PHY_3980 ();
 sky130_fd_sc_hd__decap_3 PHY_3981 ();
 sky130_fd_sc_hd__decap_3 PHY_3982 ();
 sky130_fd_sc_hd__decap_3 PHY_3983 ();
 sky130_fd_sc_hd__decap_3 PHY_3984 ();
 sky130_fd_sc_hd__decap_3 PHY_3985 ();
 sky130_fd_sc_hd__decap_3 PHY_3986 ();
 sky130_fd_sc_hd__decap_3 PHY_3987 ();
 sky130_fd_sc_hd__decap_3 PHY_3988 ();
 sky130_fd_sc_hd__decap_3 PHY_3989 ();
 sky130_fd_sc_hd__decap_3 PHY_3990 ();
 sky130_fd_sc_hd__decap_3 PHY_3991 ();
 sky130_fd_sc_hd__decap_3 PHY_3992 ();
 sky130_fd_sc_hd__decap_3 PHY_3993 ();
 sky130_fd_sc_hd__decap_3 PHY_3994 ();
 sky130_fd_sc_hd__decap_3 PHY_3995 ();
 sky130_fd_sc_hd__decap_3 PHY_3996 ();
 sky130_fd_sc_hd__decap_3 PHY_3997 ();
 sky130_fd_sc_hd__decap_3 PHY_3998 ();
 sky130_fd_sc_hd__decap_3 PHY_3999 ();
 sky130_fd_sc_hd__decap_3 PHY_4000 ();
 sky130_fd_sc_hd__decap_3 PHY_4001 ();
 sky130_fd_sc_hd__decap_3 PHY_4002 ();
 sky130_fd_sc_hd__decap_3 PHY_4003 ();
 sky130_fd_sc_hd__decap_3 PHY_4004 ();
 sky130_fd_sc_hd__decap_3 PHY_4005 ();
 sky130_fd_sc_hd__decap_3 PHY_4006 ();
 sky130_fd_sc_hd__decap_3 PHY_4007 ();
 sky130_fd_sc_hd__decap_3 PHY_4008 ();
 sky130_fd_sc_hd__decap_3 PHY_4009 ();
 sky130_fd_sc_hd__decap_3 PHY_4010 ();
 sky130_fd_sc_hd__decap_3 PHY_4011 ();
 sky130_fd_sc_hd__decap_3 PHY_4012 ();
 sky130_fd_sc_hd__decap_3 PHY_4013 ();
 sky130_fd_sc_hd__decap_3 PHY_4014 ();
 sky130_fd_sc_hd__decap_3 PHY_4015 ();
 sky130_fd_sc_hd__decap_3 PHY_4016 ();
 sky130_fd_sc_hd__decap_3 PHY_4017 ();
 sky130_fd_sc_hd__decap_3 PHY_4018 ();
 sky130_fd_sc_hd__decap_3 PHY_4019 ();
 sky130_fd_sc_hd__decap_3 PHY_4020 ();
 sky130_fd_sc_hd__decap_3 PHY_4021 ();
 sky130_fd_sc_hd__decap_3 PHY_4022 ();
 sky130_fd_sc_hd__decap_3 PHY_4023 ();
 sky130_fd_sc_hd__decap_3 PHY_4024 ();
 sky130_fd_sc_hd__decap_3 PHY_4025 ();
 sky130_fd_sc_hd__decap_3 PHY_4026 ();
 sky130_fd_sc_hd__decap_3 PHY_4027 ();
 sky130_fd_sc_hd__decap_3 PHY_4028 ();
 sky130_fd_sc_hd__decap_3 PHY_4029 ();
 sky130_fd_sc_hd__decap_3 PHY_4030 ();
 sky130_fd_sc_hd__decap_3 PHY_4031 ();
 sky130_fd_sc_hd__decap_3 PHY_4032 ();
 sky130_fd_sc_hd__decap_3 PHY_4033 ();
 sky130_fd_sc_hd__decap_3 PHY_4034 ();
 sky130_fd_sc_hd__decap_3 PHY_4035 ();
 sky130_fd_sc_hd__decap_3 PHY_4036 ();
 sky130_fd_sc_hd__decap_3 PHY_4037 ();
 sky130_fd_sc_hd__decap_3 PHY_4038 ();
 sky130_fd_sc_hd__decap_3 PHY_4039 ();
 sky130_fd_sc_hd__decap_3 PHY_4040 ();
 sky130_fd_sc_hd__decap_3 PHY_4041 ();
 sky130_fd_sc_hd__decap_3 PHY_4042 ();
 sky130_fd_sc_hd__decap_3 PHY_4043 ();
 sky130_fd_sc_hd__decap_3 PHY_4044 ();
 sky130_fd_sc_hd__decap_3 PHY_4045 ();
 sky130_fd_sc_hd__decap_3 PHY_4046 ();
 sky130_fd_sc_hd__decap_3 PHY_4047 ();
 sky130_fd_sc_hd__decap_3 PHY_4048 ();
 sky130_fd_sc_hd__decap_3 PHY_4049 ();
 sky130_fd_sc_hd__decap_3 PHY_4050 ();
 sky130_fd_sc_hd__decap_3 PHY_4051 ();
 sky130_fd_sc_hd__decap_3 PHY_4052 ();
 sky130_fd_sc_hd__decap_3 PHY_4053 ();
 sky130_fd_sc_hd__decap_3 PHY_4054 ();
 sky130_fd_sc_hd__decap_3 PHY_4055 ();
 sky130_fd_sc_hd__decap_3 PHY_4056 ();
 sky130_fd_sc_hd__decap_3 PHY_4057 ();
 sky130_fd_sc_hd__decap_3 PHY_4058 ();
 sky130_fd_sc_hd__decap_3 PHY_4059 ();
 sky130_fd_sc_hd__decap_3 PHY_4060 ();
 sky130_fd_sc_hd__decap_3 PHY_4061 ();
 sky130_fd_sc_hd__decap_3 PHY_4062 ();
 sky130_fd_sc_hd__decap_3 PHY_4063 ();
 sky130_fd_sc_hd__decap_3 PHY_4064 ();
 sky130_fd_sc_hd__decap_3 PHY_4065 ();
 sky130_fd_sc_hd__decap_3 PHY_4066 ();
 sky130_fd_sc_hd__decap_3 PHY_4067 ();
 sky130_fd_sc_hd__decap_3 PHY_4068 ();
 sky130_fd_sc_hd__decap_3 PHY_4069 ();
 sky130_fd_sc_hd__decap_3 PHY_4070 ();
 sky130_fd_sc_hd__decap_3 PHY_4071 ();
 sky130_fd_sc_hd__decap_3 PHY_4072 ();
 sky130_fd_sc_hd__decap_3 PHY_4073 ();
 sky130_fd_sc_hd__decap_3 PHY_4074 ();
 sky130_fd_sc_hd__decap_3 PHY_4075 ();
 sky130_fd_sc_hd__decap_3 PHY_4076 ();
 sky130_fd_sc_hd__decap_3 PHY_4077 ();
 sky130_fd_sc_hd__decap_3 PHY_4078 ();
 sky130_fd_sc_hd__decap_3 PHY_4079 ();
 sky130_fd_sc_hd__decap_3 PHY_4080 ();
 sky130_fd_sc_hd__decap_3 PHY_4081 ();
 sky130_fd_sc_hd__decap_3 PHY_4082 ();
 sky130_fd_sc_hd__decap_3 PHY_4083 ();
 sky130_fd_sc_hd__decap_3 PHY_4084 ();
 sky130_fd_sc_hd__decap_3 PHY_4085 ();
 sky130_fd_sc_hd__decap_3 PHY_4086 ();
 sky130_fd_sc_hd__decap_3 PHY_4087 ();
 sky130_fd_sc_hd__decap_3 PHY_4088 ();
 sky130_fd_sc_hd__decap_3 PHY_4089 ();
 sky130_fd_sc_hd__decap_3 PHY_4090 ();
 sky130_fd_sc_hd__decap_3 PHY_4091 ();
 sky130_fd_sc_hd__decap_3 PHY_4092 ();
 sky130_fd_sc_hd__decap_3 PHY_4093 ();
 sky130_fd_sc_hd__decap_3 PHY_4094 ();
 sky130_fd_sc_hd__decap_3 PHY_4095 ();
 sky130_fd_sc_hd__decap_3 PHY_4096 ();
 sky130_fd_sc_hd__decap_3 PHY_4097 ();
 sky130_fd_sc_hd__decap_3 PHY_4098 ();
 sky130_fd_sc_hd__decap_3 PHY_4099 ();
 sky130_fd_sc_hd__decap_3 PHY_4100 ();
 sky130_fd_sc_hd__decap_3 PHY_4101 ();
 sky130_fd_sc_hd__decap_3 PHY_4102 ();
 sky130_fd_sc_hd__decap_3 PHY_4103 ();
 sky130_fd_sc_hd__decap_3 PHY_4104 ();
 sky130_fd_sc_hd__decap_3 PHY_4105 ();
 sky130_fd_sc_hd__decap_3 PHY_4106 ();
 sky130_fd_sc_hd__decap_3 PHY_4107 ();
 sky130_fd_sc_hd__decap_3 PHY_4108 ();
 sky130_fd_sc_hd__decap_3 PHY_4109 ();
 sky130_fd_sc_hd__decap_3 PHY_4110 ();
 sky130_fd_sc_hd__decap_3 PHY_4111 ();
 sky130_fd_sc_hd__decap_3 PHY_4112 ();
 sky130_fd_sc_hd__decap_3 PHY_4113 ();
 sky130_fd_sc_hd__decap_3 PHY_4114 ();
 sky130_fd_sc_hd__decap_3 PHY_4115 ();
 sky130_fd_sc_hd__decap_3 PHY_4116 ();
 sky130_fd_sc_hd__decap_3 PHY_4117 ();
 sky130_fd_sc_hd__decap_3 PHY_4118 ();
 sky130_fd_sc_hd__decap_3 PHY_4119 ();
 sky130_fd_sc_hd__decap_3 PHY_4120 ();
 sky130_fd_sc_hd__decap_3 PHY_4121 ();
 sky130_fd_sc_hd__decap_3 PHY_4122 ();
 sky130_fd_sc_hd__decap_3 PHY_4123 ();
 sky130_fd_sc_hd__decap_3 PHY_4124 ();
 sky130_fd_sc_hd__decap_3 PHY_4125 ();
 sky130_fd_sc_hd__decap_3 PHY_4126 ();
 sky130_fd_sc_hd__decap_3 PHY_4127 ();
 sky130_fd_sc_hd__decap_3 PHY_4128 ();
 sky130_fd_sc_hd__decap_3 PHY_4129 ();
 sky130_fd_sc_hd__decap_3 PHY_4130 ();
 sky130_fd_sc_hd__decap_3 PHY_4131 ();
 sky130_fd_sc_hd__decap_3 PHY_4132 ();
 sky130_fd_sc_hd__decap_3 PHY_4133 ();
 sky130_fd_sc_hd__decap_3 PHY_4134 ();
 sky130_fd_sc_hd__decap_3 PHY_4135 ();
 sky130_fd_sc_hd__decap_3 PHY_4136 ();
 sky130_fd_sc_hd__decap_3 PHY_4137 ();
 sky130_fd_sc_hd__decap_3 PHY_4138 ();
 sky130_fd_sc_hd__decap_3 PHY_4139 ();
 sky130_fd_sc_hd__decap_3 PHY_4140 ();
 sky130_fd_sc_hd__decap_3 PHY_4141 ();
 sky130_fd_sc_hd__decap_3 PHY_4142 ();
 sky130_fd_sc_hd__decap_3 PHY_4143 ();
 sky130_fd_sc_hd__decap_3 PHY_4144 ();
 sky130_fd_sc_hd__decap_3 PHY_4145 ();
 sky130_fd_sc_hd__decap_3 PHY_4146 ();
 sky130_fd_sc_hd__decap_3 PHY_4147 ();
 sky130_fd_sc_hd__decap_3 PHY_4148 ();
 sky130_fd_sc_hd__decap_3 PHY_4149 ();
 sky130_fd_sc_hd__decap_3 PHY_4150 ();
 sky130_fd_sc_hd__decap_3 PHY_4151 ();
 sky130_fd_sc_hd__decap_3 PHY_4152 ();
 sky130_fd_sc_hd__decap_3 PHY_4153 ();
 sky130_fd_sc_hd__decap_3 PHY_4154 ();
 sky130_fd_sc_hd__decap_3 PHY_4155 ();
 sky130_fd_sc_hd__decap_3 PHY_4156 ();
 sky130_fd_sc_hd__decap_3 PHY_4157 ();
 sky130_fd_sc_hd__decap_3 PHY_4158 ();
 sky130_fd_sc_hd__decap_3 PHY_4159 ();
 sky130_fd_sc_hd__decap_3 PHY_4160 ();
 sky130_fd_sc_hd__decap_3 PHY_4161 ();
 sky130_fd_sc_hd__decap_3 PHY_4162 ();
 sky130_fd_sc_hd__decap_3 PHY_4163 ();
 sky130_fd_sc_hd__decap_3 PHY_4164 ();
 sky130_fd_sc_hd__decap_3 PHY_4165 ();
 sky130_fd_sc_hd__decap_3 PHY_4166 ();
 sky130_fd_sc_hd__decap_3 PHY_4167 ();
 sky130_fd_sc_hd__decap_3 PHY_4168 ();
 sky130_fd_sc_hd__decap_3 PHY_4169 ();
 sky130_fd_sc_hd__decap_3 PHY_4170 ();
 sky130_fd_sc_hd__decap_3 PHY_4171 ();
 sky130_fd_sc_hd__decap_3 PHY_4172 ();
 sky130_fd_sc_hd__decap_3 PHY_4173 ();
 sky130_fd_sc_hd__decap_3 PHY_4174 ();
 sky130_fd_sc_hd__decap_3 PHY_4175 ();
 sky130_fd_sc_hd__decap_3 PHY_4176 ();
 sky130_fd_sc_hd__decap_3 PHY_4177 ();
 sky130_fd_sc_hd__decap_3 PHY_4178 ();
 sky130_fd_sc_hd__decap_3 PHY_4179 ();
 sky130_fd_sc_hd__decap_3 PHY_4180 ();
 sky130_fd_sc_hd__decap_3 PHY_4181 ();
 sky130_fd_sc_hd__decap_3 PHY_4182 ();
 sky130_fd_sc_hd__decap_3 PHY_4183 ();
 sky130_fd_sc_hd__decap_3 PHY_4184 ();
 sky130_fd_sc_hd__decap_3 PHY_4185 ();
 sky130_fd_sc_hd__decap_3 PHY_4186 ();
 sky130_fd_sc_hd__decap_3 PHY_4187 ();
 sky130_fd_sc_hd__decap_3 PHY_4188 ();
 sky130_fd_sc_hd__decap_3 PHY_4189 ();
 sky130_fd_sc_hd__decap_3 PHY_4190 ();
 sky130_fd_sc_hd__decap_3 PHY_4191 ();
 sky130_fd_sc_hd__decap_3 PHY_4192 ();
 sky130_fd_sc_hd__decap_3 PHY_4193 ();
 sky130_fd_sc_hd__decap_3 PHY_4194 ();
 sky130_fd_sc_hd__decap_3 PHY_4195 ();
 sky130_fd_sc_hd__decap_3 PHY_4196 ();
 sky130_fd_sc_hd__decap_3 PHY_4197 ();
 sky130_fd_sc_hd__decap_3 PHY_4198 ();
 sky130_fd_sc_hd__decap_3 PHY_4199 ();
 sky130_fd_sc_hd__decap_3 PHY_4200 ();
 sky130_fd_sc_hd__decap_3 PHY_4201 ();
 sky130_fd_sc_hd__decap_3 PHY_4202 ();
 sky130_fd_sc_hd__decap_3 PHY_4203 ();
 sky130_fd_sc_hd__decap_3 PHY_4204 ();
 sky130_fd_sc_hd__decap_3 PHY_4205 ();
 sky130_fd_sc_hd__decap_3 PHY_4206 ();
 sky130_fd_sc_hd__decap_3 PHY_4207 ();
 sky130_fd_sc_hd__decap_3 PHY_4208 ();
 sky130_fd_sc_hd__decap_3 PHY_4209 ();
 sky130_fd_sc_hd__decap_3 PHY_4210 ();
 sky130_fd_sc_hd__decap_3 PHY_4211 ();
 sky130_fd_sc_hd__decap_3 PHY_4212 ();
 sky130_fd_sc_hd__decap_3 PHY_4213 ();
 sky130_fd_sc_hd__decap_3 PHY_4214 ();
 sky130_fd_sc_hd__decap_3 PHY_4215 ();
 sky130_fd_sc_hd__decap_3 PHY_4216 ();
 sky130_fd_sc_hd__decap_3 PHY_4217 ();
 sky130_fd_sc_hd__decap_3 PHY_4218 ();
 sky130_fd_sc_hd__decap_3 PHY_4219 ();
 sky130_fd_sc_hd__decap_3 PHY_4220 ();
 sky130_fd_sc_hd__decap_3 PHY_4221 ();
 sky130_fd_sc_hd__decap_3 PHY_4222 ();
 sky130_fd_sc_hd__decap_3 PHY_4223 ();
 sky130_fd_sc_hd__decap_3 PHY_4224 ();
 sky130_fd_sc_hd__decap_3 PHY_4225 ();
 sky130_fd_sc_hd__decap_3 PHY_4226 ();
 sky130_fd_sc_hd__decap_3 PHY_4227 ();
 sky130_fd_sc_hd__decap_3 PHY_4228 ();
 sky130_fd_sc_hd__decap_3 PHY_4229 ();
 sky130_fd_sc_hd__decap_3 PHY_4230 ();
 sky130_fd_sc_hd__decap_3 PHY_4231 ();
 sky130_fd_sc_hd__decap_3 PHY_4232 ();
 sky130_fd_sc_hd__decap_3 PHY_4233 ();
 sky130_fd_sc_hd__decap_3 PHY_4234 ();
 sky130_fd_sc_hd__decap_3 PHY_4235 ();
 sky130_fd_sc_hd__decap_3 PHY_4236 ();
 sky130_fd_sc_hd__decap_3 PHY_4237 ();
 sky130_fd_sc_hd__decap_3 PHY_4238 ();
 sky130_fd_sc_hd__decap_3 PHY_4239 ();
 sky130_fd_sc_hd__decap_3 PHY_4240 ();
 sky130_fd_sc_hd__decap_3 PHY_4241 ();
 sky130_fd_sc_hd__decap_3 PHY_4242 ();
 sky130_fd_sc_hd__decap_3 PHY_4243 ();
 sky130_fd_sc_hd__decap_3 PHY_4244 ();
 sky130_fd_sc_hd__decap_3 PHY_4245 ();
 sky130_fd_sc_hd__decap_3 PHY_4246 ();
 sky130_fd_sc_hd__decap_3 PHY_4247 ();
 sky130_fd_sc_hd__decap_3 PHY_4248 ();
 sky130_fd_sc_hd__decap_3 PHY_4249 ();
 sky130_fd_sc_hd__decap_3 PHY_4250 ();
 sky130_fd_sc_hd__decap_3 PHY_4251 ();
 sky130_fd_sc_hd__decap_3 PHY_4252 ();
 sky130_fd_sc_hd__decap_3 PHY_4253 ();
 sky130_fd_sc_hd__decap_3 PHY_4254 ();
 sky130_fd_sc_hd__decap_3 PHY_4255 ();
 sky130_fd_sc_hd__decap_3 PHY_4256 ();
 sky130_fd_sc_hd__decap_3 PHY_4257 ();
 sky130_fd_sc_hd__decap_3 PHY_4258 ();
 sky130_fd_sc_hd__decap_3 PHY_4259 ();
 sky130_fd_sc_hd__decap_3 PHY_4260 ();
 sky130_fd_sc_hd__decap_3 PHY_4261 ();
 sky130_fd_sc_hd__decap_3 PHY_4262 ();
 sky130_fd_sc_hd__decap_3 PHY_4263 ();
 sky130_fd_sc_hd__decap_3 PHY_4264 ();
 sky130_fd_sc_hd__decap_3 PHY_4265 ();
 sky130_fd_sc_hd__decap_3 PHY_4266 ();
 sky130_fd_sc_hd__decap_3 PHY_4267 ();
 sky130_fd_sc_hd__decap_3 PHY_4268 ();
 sky130_fd_sc_hd__decap_3 PHY_4269 ();
 sky130_fd_sc_hd__decap_3 PHY_4270 ();
 sky130_fd_sc_hd__decap_3 PHY_4271 ();
 sky130_fd_sc_hd__decap_3 PHY_4272 ();
 sky130_fd_sc_hd__decap_3 PHY_4273 ();
 sky130_fd_sc_hd__decap_3 PHY_4274 ();
 sky130_fd_sc_hd__decap_3 PHY_4275 ();
 sky130_fd_sc_hd__decap_3 PHY_4276 ();
 sky130_fd_sc_hd__decap_3 PHY_4277 ();
 sky130_fd_sc_hd__decap_3 PHY_4278 ();
 sky130_fd_sc_hd__decap_3 PHY_4279 ();
 sky130_fd_sc_hd__decap_3 PHY_4280 ();
 sky130_fd_sc_hd__decap_3 PHY_4281 ();
 sky130_fd_sc_hd__decap_3 PHY_4282 ();
 sky130_fd_sc_hd__decap_3 PHY_4283 ();
 sky130_fd_sc_hd__decap_3 PHY_4284 ();
 sky130_fd_sc_hd__decap_3 PHY_4285 ();
 sky130_fd_sc_hd__decap_3 PHY_4286 ();
 sky130_fd_sc_hd__decap_3 PHY_4287 ();
 sky130_fd_sc_hd__decap_3 PHY_4288 ();
 sky130_fd_sc_hd__decap_3 PHY_4289 ();
 sky130_fd_sc_hd__decap_3 PHY_4290 ();
 sky130_fd_sc_hd__decap_3 PHY_4291 ();
 sky130_fd_sc_hd__decap_3 PHY_4292 ();
 sky130_fd_sc_hd__decap_3 PHY_4293 ();
 sky130_fd_sc_hd__decap_3 PHY_4294 ();
 sky130_fd_sc_hd__decap_3 PHY_4295 ();
 sky130_fd_sc_hd__decap_3 PHY_4296 ();
 sky130_fd_sc_hd__decap_3 PHY_4297 ();
 sky130_fd_sc_hd__decap_3 PHY_4298 ();
 sky130_fd_sc_hd__decap_3 PHY_4299 ();
 sky130_fd_sc_hd__decap_3 PHY_4300 ();
 sky130_fd_sc_hd__decap_3 PHY_4301 ();
 sky130_fd_sc_hd__decap_3 PHY_4302 ();
 sky130_fd_sc_hd__decap_3 PHY_4303 ();
 sky130_fd_sc_hd__decap_3 PHY_4304 ();
 sky130_fd_sc_hd__decap_3 PHY_4305 ();
 sky130_fd_sc_hd__decap_3 PHY_4306 ();
 sky130_fd_sc_hd__decap_3 PHY_4307 ();
 sky130_fd_sc_hd__decap_3 PHY_4308 ();
 sky130_fd_sc_hd__decap_3 PHY_4309 ();
 sky130_fd_sc_hd__decap_3 PHY_4310 ();
 sky130_fd_sc_hd__decap_3 PHY_4311 ();
 sky130_fd_sc_hd__decap_3 PHY_4312 ();
 sky130_fd_sc_hd__decap_3 PHY_4313 ();
 sky130_fd_sc_hd__decap_3 PHY_4314 ();
 sky130_fd_sc_hd__decap_3 PHY_4315 ();
 sky130_fd_sc_hd__decap_3 PHY_4316 ();
 sky130_fd_sc_hd__decap_3 PHY_4317 ();
 sky130_fd_sc_hd__decap_3 PHY_4318 ();
 sky130_fd_sc_hd__decap_3 PHY_4319 ();
 sky130_fd_sc_hd__decap_3 PHY_4320 ();
 sky130_fd_sc_hd__decap_3 PHY_4321 ();
 sky130_fd_sc_hd__decap_3 PHY_4322 ();
 sky130_fd_sc_hd__decap_3 PHY_4323 ();
 sky130_fd_sc_hd__decap_3 PHY_4324 ();
 sky130_fd_sc_hd__decap_3 PHY_4325 ();
 sky130_fd_sc_hd__decap_3 PHY_4326 ();
 sky130_fd_sc_hd__decap_3 PHY_4327 ();
 sky130_fd_sc_hd__decap_3 PHY_4328 ();
 sky130_fd_sc_hd__decap_3 PHY_4329 ();
 sky130_fd_sc_hd__decap_3 PHY_4330 ();
 sky130_fd_sc_hd__decap_3 PHY_4331 ();
 sky130_fd_sc_hd__decap_3 PHY_4332 ();
 sky130_fd_sc_hd__decap_3 PHY_4333 ();
 sky130_fd_sc_hd__decap_3 PHY_4334 ();
 sky130_fd_sc_hd__decap_3 PHY_4335 ();
 sky130_fd_sc_hd__decap_3 PHY_4336 ();
 sky130_fd_sc_hd__decap_3 PHY_4337 ();
 sky130_fd_sc_hd__decap_3 PHY_4338 ();
 sky130_fd_sc_hd__decap_3 PHY_4339 ();
 sky130_fd_sc_hd__decap_3 PHY_4340 ();
 sky130_fd_sc_hd__decap_3 PHY_4341 ();
 sky130_fd_sc_hd__decap_3 PHY_4342 ();
 sky130_fd_sc_hd__decap_3 PHY_4343 ();
 sky130_fd_sc_hd__decap_3 PHY_4344 ();
 sky130_fd_sc_hd__decap_3 PHY_4345 ();
 sky130_fd_sc_hd__decap_3 PHY_4346 ();
 sky130_fd_sc_hd__decap_3 PHY_4347 ();
 sky130_fd_sc_hd__decap_3 PHY_4348 ();
 sky130_fd_sc_hd__decap_3 PHY_4349 ();
 sky130_fd_sc_hd__decap_3 PHY_4350 ();
 sky130_fd_sc_hd__decap_3 PHY_4351 ();
 sky130_fd_sc_hd__decap_3 PHY_4352 ();
 sky130_fd_sc_hd__decap_3 PHY_4353 ();
 sky130_fd_sc_hd__decap_3 PHY_4354 ();
 sky130_fd_sc_hd__decap_3 PHY_4355 ();
 sky130_fd_sc_hd__decap_3 PHY_4356 ();
 sky130_fd_sc_hd__decap_3 PHY_4357 ();
 sky130_fd_sc_hd__decap_3 PHY_4358 ();
 sky130_fd_sc_hd__decap_3 PHY_4359 ();
 sky130_fd_sc_hd__decap_3 PHY_4360 ();
 sky130_fd_sc_hd__decap_3 PHY_4361 ();
 sky130_fd_sc_hd__decap_3 PHY_4362 ();
 sky130_fd_sc_hd__decap_3 PHY_4363 ();
 sky130_fd_sc_hd__decap_3 PHY_4364 ();
 sky130_fd_sc_hd__decap_3 PHY_4365 ();
 sky130_fd_sc_hd__decap_3 PHY_4366 ();
 sky130_fd_sc_hd__decap_3 PHY_4367 ();
 sky130_fd_sc_hd__decap_3 PHY_4368 ();
 sky130_fd_sc_hd__decap_3 PHY_4369 ();
 sky130_fd_sc_hd__decap_3 PHY_4370 ();
 sky130_fd_sc_hd__decap_3 PHY_4371 ();
 sky130_fd_sc_hd__decap_3 PHY_4372 ();
 sky130_fd_sc_hd__decap_3 PHY_4373 ();
 sky130_fd_sc_hd__decap_3 PHY_4374 ();
 sky130_fd_sc_hd__decap_3 PHY_4375 ();
 sky130_fd_sc_hd__decap_3 PHY_4376 ();
 sky130_fd_sc_hd__decap_3 PHY_4377 ();
 sky130_fd_sc_hd__decap_3 PHY_4378 ();
 sky130_fd_sc_hd__decap_3 PHY_4379 ();
 sky130_fd_sc_hd__decap_3 PHY_4380 ();
 sky130_fd_sc_hd__decap_3 PHY_4381 ();
 sky130_fd_sc_hd__decap_3 PHY_4382 ();
 sky130_fd_sc_hd__decap_3 PHY_4383 ();
 sky130_fd_sc_hd__decap_3 PHY_4384 ();
 sky130_fd_sc_hd__decap_3 PHY_4385 ();
 sky130_fd_sc_hd__decap_3 PHY_4386 ();
 sky130_fd_sc_hd__decap_3 PHY_4387 ();
 sky130_fd_sc_hd__decap_3 PHY_4388 ();
 sky130_fd_sc_hd__decap_3 PHY_4389 ();
 sky130_fd_sc_hd__decap_3 PHY_4390 ();
 sky130_fd_sc_hd__decap_3 PHY_4391 ();
 sky130_fd_sc_hd__decap_3 PHY_4392 ();
 sky130_fd_sc_hd__decap_3 PHY_4393 ();
 sky130_fd_sc_hd__decap_3 PHY_4394 ();
 sky130_fd_sc_hd__decap_3 PHY_4395 ();
 sky130_fd_sc_hd__decap_3 PHY_4396 ();
 sky130_fd_sc_hd__decap_3 PHY_4397 ();
 sky130_fd_sc_hd__decap_3 PHY_4398 ();
 sky130_fd_sc_hd__decap_3 PHY_4399 ();
 sky130_fd_sc_hd__decap_3 PHY_4400 ();
 sky130_fd_sc_hd__decap_3 PHY_4401 ();
 sky130_fd_sc_hd__decap_3 PHY_4402 ();
 sky130_fd_sc_hd__decap_3 PHY_4403 ();
 sky130_fd_sc_hd__decap_3 PHY_4404 ();
 sky130_fd_sc_hd__decap_3 PHY_4405 ();
 sky130_fd_sc_hd__decap_3 PHY_4406 ();
 sky130_fd_sc_hd__decap_3 PHY_4407 ();
 sky130_fd_sc_hd__decap_3 PHY_4408 ();
 sky130_fd_sc_hd__decap_3 PHY_4409 ();
 sky130_fd_sc_hd__decap_3 PHY_4410 ();
 sky130_fd_sc_hd__decap_3 PHY_4411 ();
 sky130_fd_sc_hd__decap_3 PHY_4412 ();
 sky130_fd_sc_hd__decap_3 PHY_4413 ();
 sky130_fd_sc_hd__decap_3 PHY_4414 ();
 sky130_fd_sc_hd__decap_3 PHY_4415 ();
 sky130_fd_sc_hd__decap_3 PHY_4416 ();
 sky130_fd_sc_hd__decap_3 PHY_4417 ();
 sky130_fd_sc_hd__decap_3 PHY_4418 ();
 sky130_fd_sc_hd__decap_3 PHY_4419 ();
 sky130_fd_sc_hd__decap_3 PHY_4420 ();
 sky130_fd_sc_hd__decap_3 PHY_4421 ();
 sky130_fd_sc_hd__decap_3 PHY_4422 ();
 sky130_fd_sc_hd__decap_3 PHY_4423 ();
 sky130_fd_sc_hd__decap_3 PHY_4424 ();
 sky130_fd_sc_hd__decap_3 PHY_4425 ();
 sky130_fd_sc_hd__decap_3 PHY_4426 ();
 sky130_fd_sc_hd__decap_3 PHY_4427 ();
 sky130_fd_sc_hd__decap_3 PHY_4428 ();
 sky130_fd_sc_hd__decap_3 PHY_4429 ();
 sky130_fd_sc_hd__decap_3 PHY_4430 ();
 sky130_fd_sc_hd__decap_3 PHY_4431 ();
 sky130_fd_sc_hd__decap_3 PHY_4432 ();
 sky130_fd_sc_hd__decap_3 PHY_4433 ();
 sky130_fd_sc_hd__decap_3 PHY_4434 ();
 sky130_fd_sc_hd__decap_3 PHY_4435 ();
 sky130_fd_sc_hd__decap_3 PHY_4436 ();
 sky130_fd_sc_hd__decap_3 PHY_4437 ();
 sky130_fd_sc_hd__decap_3 PHY_4438 ();
 sky130_fd_sc_hd__decap_3 PHY_4439 ();
 sky130_fd_sc_hd__decap_3 PHY_4440 ();
 sky130_fd_sc_hd__decap_3 PHY_4441 ();
 sky130_fd_sc_hd__decap_3 PHY_4442 ();
 sky130_fd_sc_hd__decap_3 PHY_4443 ();
 sky130_fd_sc_hd__decap_3 PHY_4444 ();
 sky130_fd_sc_hd__decap_3 PHY_4445 ();
 sky130_fd_sc_hd__decap_3 PHY_4446 ();
 sky130_fd_sc_hd__decap_3 PHY_4447 ();
 sky130_fd_sc_hd__decap_3 PHY_4448 ();
 sky130_fd_sc_hd__decap_3 PHY_4449 ();
 sky130_fd_sc_hd__decap_3 PHY_4450 ();
 sky130_fd_sc_hd__decap_3 PHY_4451 ();
 sky130_fd_sc_hd__decap_3 PHY_4452 ();
 sky130_fd_sc_hd__decap_3 PHY_4453 ();
 sky130_fd_sc_hd__decap_3 PHY_4454 ();
 sky130_fd_sc_hd__decap_3 PHY_4455 ();
 sky130_fd_sc_hd__decap_3 PHY_4456 ();
 sky130_fd_sc_hd__decap_3 PHY_4457 ();
 sky130_fd_sc_hd__decap_3 PHY_4458 ();
 sky130_fd_sc_hd__decap_3 PHY_4459 ();
 sky130_fd_sc_hd__decap_3 PHY_4460 ();
 sky130_fd_sc_hd__decap_3 PHY_4461 ();
 sky130_fd_sc_hd__decap_3 PHY_4462 ();
 sky130_fd_sc_hd__decap_3 PHY_4463 ();
 sky130_fd_sc_hd__decap_3 PHY_4464 ();
 sky130_fd_sc_hd__decap_3 PHY_4465 ();
 sky130_fd_sc_hd__decap_3 PHY_4466 ();
 sky130_fd_sc_hd__decap_3 PHY_4467 ();
 sky130_fd_sc_hd__decap_3 PHY_4468 ();
 sky130_fd_sc_hd__decap_3 PHY_4469 ();
 sky130_fd_sc_hd__decap_3 PHY_4470 ();
 sky130_fd_sc_hd__decap_3 PHY_4471 ();
 sky130_fd_sc_hd__decap_3 PHY_4472 ();
 sky130_fd_sc_hd__decap_3 PHY_4473 ();
 sky130_fd_sc_hd__decap_3 PHY_4474 ();
 sky130_fd_sc_hd__decap_3 PHY_4475 ();
 sky130_fd_sc_hd__decap_3 PHY_4476 ();
 sky130_fd_sc_hd__decap_3 PHY_4477 ();
 sky130_fd_sc_hd__decap_3 PHY_4478 ();
 sky130_fd_sc_hd__decap_3 PHY_4479 ();
 sky130_fd_sc_hd__decap_3 PHY_4480 ();
 sky130_fd_sc_hd__decap_3 PHY_4481 ();
 sky130_fd_sc_hd__decap_3 PHY_4482 ();
 sky130_fd_sc_hd__decap_3 PHY_4483 ();
 sky130_fd_sc_hd__decap_3 PHY_4484 ();
 sky130_fd_sc_hd__decap_3 PHY_4485 ();
 sky130_fd_sc_hd__decap_3 PHY_4486 ();
 sky130_fd_sc_hd__decap_3 PHY_4487 ();
 sky130_fd_sc_hd__decap_3 PHY_4488 ();
 sky130_fd_sc_hd__decap_3 PHY_4489 ();
 sky130_fd_sc_hd__decap_3 PHY_4490 ();
 sky130_fd_sc_hd__decap_3 PHY_4491 ();
 sky130_fd_sc_hd__decap_3 PHY_4492 ();
 sky130_fd_sc_hd__decap_3 PHY_4493 ();
 sky130_fd_sc_hd__decap_3 PHY_4494 ();
 sky130_fd_sc_hd__decap_3 PHY_4495 ();
 sky130_fd_sc_hd__decap_3 PHY_4496 ();
 sky130_fd_sc_hd__decap_3 PHY_4497 ();
 sky130_fd_sc_hd__decap_3 PHY_4498 ();
 sky130_fd_sc_hd__decap_3 PHY_4499 ();
 sky130_fd_sc_hd__decap_3 PHY_4500 ();
 sky130_fd_sc_hd__decap_3 PHY_4501 ();
 sky130_fd_sc_hd__decap_3 PHY_4502 ();
 sky130_fd_sc_hd__decap_3 PHY_4503 ();
 sky130_fd_sc_hd__decap_3 PHY_4504 ();
 sky130_fd_sc_hd__decap_3 PHY_4505 ();
 sky130_fd_sc_hd__decap_3 PHY_4506 ();
 sky130_fd_sc_hd__decap_3 PHY_4507 ();
 sky130_fd_sc_hd__decap_3 PHY_4508 ();
 sky130_fd_sc_hd__decap_3 PHY_4509 ();
 sky130_fd_sc_hd__decap_3 PHY_4510 ();
 sky130_fd_sc_hd__decap_3 PHY_4511 ();
 sky130_fd_sc_hd__decap_3 PHY_4512 ();
 sky130_fd_sc_hd__decap_3 PHY_4513 ();
 sky130_fd_sc_hd__decap_3 PHY_4514 ();
 sky130_fd_sc_hd__decap_3 PHY_4515 ();
 sky130_fd_sc_hd__decap_3 PHY_4516 ();
 sky130_fd_sc_hd__decap_3 PHY_4517 ();
 sky130_fd_sc_hd__decap_3 PHY_4518 ();
 sky130_fd_sc_hd__decap_3 PHY_4519 ();
 sky130_fd_sc_hd__decap_3 PHY_4520 ();
 sky130_fd_sc_hd__decap_3 PHY_4521 ();
 sky130_fd_sc_hd__decap_3 PHY_4522 ();
 sky130_fd_sc_hd__decap_3 PHY_4523 ();
 sky130_fd_sc_hd__decap_3 PHY_4524 ();
 sky130_fd_sc_hd__decap_3 PHY_4525 ();
 sky130_fd_sc_hd__decap_3 PHY_4526 ();
 sky130_fd_sc_hd__decap_3 PHY_4527 ();
 sky130_fd_sc_hd__decap_3 PHY_4528 ();
 sky130_fd_sc_hd__decap_3 PHY_4529 ();
 sky130_fd_sc_hd__decap_3 PHY_4530 ();
 sky130_fd_sc_hd__decap_3 PHY_4531 ();
 sky130_fd_sc_hd__decap_3 PHY_4532 ();
 sky130_fd_sc_hd__decap_3 PHY_4533 ();
 sky130_fd_sc_hd__decap_3 PHY_4534 ();
 sky130_fd_sc_hd__decap_3 PHY_4535 ();
 sky130_fd_sc_hd__decap_3 PHY_4536 ();
 sky130_fd_sc_hd__decap_3 PHY_4537 ();
 sky130_fd_sc_hd__decap_3 PHY_4538 ();
 sky130_fd_sc_hd__decap_3 PHY_4539 ();
 sky130_fd_sc_hd__decap_3 PHY_4540 ();
 sky130_fd_sc_hd__decap_3 PHY_4541 ();
 sky130_fd_sc_hd__decap_3 PHY_4542 ();
 sky130_fd_sc_hd__decap_3 PHY_4543 ();
 sky130_fd_sc_hd__decap_3 PHY_4544 ();
 sky130_fd_sc_hd__decap_3 PHY_4545 ();
 sky130_fd_sc_hd__decap_3 PHY_4546 ();
 sky130_fd_sc_hd__decap_3 PHY_4547 ();
 sky130_fd_sc_hd__decap_3 PHY_4548 ();
 sky130_fd_sc_hd__decap_3 PHY_4549 ();
 sky130_fd_sc_hd__decap_3 PHY_4550 ();
 sky130_fd_sc_hd__decap_3 PHY_4551 ();
 sky130_fd_sc_hd__decap_3 PHY_4552 ();
 sky130_fd_sc_hd__decap_3 PHY_4553 ();
 sky130_fd_sc_hd__decap_3 PHY_4554 ();
 sky130_fd_sc_hd__decap_3 PHY_4555 ();
 sky130_fd_sc_hd__decap_3 PHY_4556 ();
 sky130_fd_sc_hd__decap_3 PHY_4557 ();
 sky130_fd_sc_hd__decap_3 PHY_4558 ();
 sky130_fd_sc_hd__decap_3 PHY_4559 ();
 sky130_fd_sc_hd__decap_3 PHY_4560 ();
 sky130_fd_sc_hd__decap_3 PHY_4561 ();
 sky130_fd_sc_hd__decap_3 PHY_4562 ();
 sky130_fd_sc_hd__decap_3 PHY_4563 ();
 sky130_fd_sc_hd__decap_3 PHY_4564 ();
 sky130_fd_sc_hd__decap_3 PHY_4565 ();
 sky130_fd_sc_hd__decap_3 PHY_4566 ();
 sky130_fd_sc_hd__decap_3 PHY_4567 ();
 sky130_fd_sc_hd__decap_3 PHY_4568 ();
 sky130_fd_sc_hd__decap_3 PHY_4569 ();
 sky130_fd_sc_hd__decap_3 PHY_4570 ();
 sky130_fd_sc_hd__decap_3 PHY_4571 ();
 sky130_fd_sc_hd__decap_3 PHY_4572 ();
 sky130_fd_sc_hd__decap_3 PHY_4573 ();
 sky130_fd_sc_hd__decap_3 PHY_4574 ();
 sky130_fd_sc_hd__decap_3 PHY_4575 ();
 sky130_fd_sc_hd__decap_3 PHY_4576 ();
 sky130_fd_sc_hd__decap_3 PHY_4577 ();
 sky130_fd_sc_hd__decap_3 PHY_4578 ();
 sky130_fd_sc_hd__decap_3 PHY_4579 ();
 sky130_fd_sc_hd__decap_3 PHY_4580 ();
 sky130_fd_sc_hd__decap_3 PHY_4581 ();
 sky130_fd_sc_hd__decap_3 PHY_4582 ();
 sky130_fd_sc_hd__decap_3 PHY_4583 ();
 sky130_fd_sc_hd__decap_3 PHY_4584 ();
 sky130_fd_sc_hd__decap_3 PHY_4585 ();
 sky130_fd_sc_hd__decap_3 PHY_4586 ();
 sky130_fd_sc_hd__decap_3 PHY_4587 ();
 sky130_fd_sc_hd__decap_3 PHY_4588 ();
 sky130_fd_sc_hd__decap_3 PHY_4589 ();
 sky130_fd_sc_hd__decap_3 PHY_4590 ();
 sky130_fd_sc_hd__decap_3 PHY_4591 ();
 sky130_fd_sc_hd__decap_3 PHY_4592 ();
 sky130_fd_sc_hd__decap_3 PHY_4593 ();
 sky130_fd_sc_hd__decap_3 PHY_4594 ();
 sky130_fd_sc_hd__decap_3 PHY_4595 ();
 sky130_fd_sc_hd__decap_3 PHY_4596 ();
 sky130_fd_sc_hd__decap_3 PHY_4597 ();
 sky130_fd_sc_hd__decap_3 PHY_4598 ();
 sky130_fd_sc_hd__decap_3 PHY_4599 ();
 sky130_fd_sc_hd__decap_3 PHY_4600 ();
 sky130_fd_sc_hd__decap_3 PHY_4601 ();
 sky130_fd_sc_hd__decap_3 PHY_4602 ();
 sky130_fd_sc_hd__decap_3 PHY_4603 ();
 sky130_fd_sc_hd__decap_3 PHY_4604 ();
 sky130_fd_sc_hd__decap_3 PHY_4605 ();
 sky130_fd_sc_hd__decap_3 PHY_4606 ();
 sky130_fd_sc_hd__decap_3 PHY_4607 ();
 sky130_fd_sc_hd__decap_3 PHY_4608 ();
 sky130_fd_sc_hd__decap_3 PHY_4609 ();
 sky130_fd_sc_hd__decap_3 PHY_4610 ();
 sky130_fd_sc_hd__decap_3 PHY_4611 ();
 sky130_fd_sc_hd__decap_3 PHY_4612 ();
 sky130_fd_sc_hd__decap_3 PHY_4613 ();
 sky130_fd_sc_hd__decap_3 PHY_4614 ();
 sky130_fd_sc_hd__decap_3 PHY_4615 ();
 sky130_fd_sc_hd__decap_3 PHY_4616 ();
 sky130_fd_sc_hd__decap_3 PHY_4617 ();
 sky130_fd_sc_hd__decap_3 PHY_4618 ();
 sky130_fd_sc_hd__decap_3 PHY_4619 ();
 sky130_fd_sc_hd__decap_3 PHY_4620 ();
 sky130_fd_sc_hd__decap_3 PHY_4621 ();
 sky130_fd_sc_hd__decap_3 PHY_4622 ();
 sky130_fd_sc_hd__decap_3 PHY_4623 ();
 sky130_fd_sc_hd__decap_3 PHY_4624 ();
 sky130_fd_sc_hd__decap_3 PHY_4625 ();
 sky130_fd_sc_hd__decap_3 PHY_4626 ();
 sky130_fd_sc_hd__decap_3 PHY_4627 ();
 sky130_fd_sc_hd__decap_3 PHY_4628 ();
 sky130_fd_sc_hd__decap_3 PHY_4629 ();
 sky130_fd_sc_hd__decap_3 PHY_4630 ();
 sky130_fd_sc_hd__decap_3 PHY_4631 ();
 sky130_fd_sc_hd__decap_3 PHY_4632 ();
 sky130_fd_sc_hd__decap_3 PHY_4633 ();
 sky130_fd_sc_hd__decap_3 PHY_4634 ();
 sky130_fd_sc_hd__decap_3 PHY_4635 ();
 sky130_fd_sc_hd__decap_3 PHY_4636 ();
 sky130_fd_sc_hd__decap_3 PHY_4637 ();
 sky130_fd_sc_hd__decap_3 PHY_4638 ();
 sky130_fd_sc_hd__decap_3 PHY_4639 ();
 sky130_fd_sc_hd__decap_3 PHY_4640 ();
 sky130_fd_sc_hd__decap_3 PHY_4641 ();
 sky130_fd_sc_hd__decap_3 PHY_4642 ();
 sky130_fd_sc_hd__decap_3 PHY_4643 ();
 sky130_fd_sc_hd__decap_3 PHY_4644 ();
 sky130_fd_sc_hd__decap_3 PHY_4645 ();
 sky130_fd_sc_hd__decap_3 PHY_4646 ();
 sky130_fd_sc_hd__decap_3 PHY_4647 ();
 sky130_fd_sc_hd__decap_3 PHY_4648 ();
 sky130_fd_sc_hd__decap_3 PHY_4649 ();
 sky130_fd_sc_hd__decap_3 PHY_4650 ();
 sky130_fd_sc_hd__decap_3 PHY_4651 ();
 sky130_fd_sc_hd__decap_3 PHY_4652 ();
 sky130_fd_sc_hd__decap_3 PHY_4653 ();
 sky130_fd_sc_hd__decap_3 PHY_4654 ();
 sky130_fd_sc_hd__decap_3 PHY_4655 ();
 sky130_fd_sc_hd__decap_3 PHY_4656 ();
 sky130_fd_sc_hd__decap_3 PHY_4657 ();
 sky130_fd_sc_hd__decap_3 PHY_4658 ();
 sky130_fd_sc_hd__decap_3 PHY_4659 ();
 sky130_fd_sc_hd__decap_3 PHY_4660 ();
 sky130_fd_sc_hd__decap_3 PHY_4661 ();
 sky130_fd_sc_hd__decap_3 PHY_4662 ();
 sky130_fd_sc_hd__decap_3 PHY_4663 ();
 sky130_fd_sc_hd__decap_3 PHY_4664 ();
 sky130_fd_sc_hd__decap_3 PHY_4665 ();
 sky130_fd_sc_hd__decap_3 PHY_4666 ();
 sky130_fd_sc_hd__decap_3 PHY_4667 ();
 sky130_fd_sc_hd__decap_3 PHY_4668 ();
 sky130_fd_sc_hd__decap_3 PHY_4669 ();
 sky130_fd_sc_hd__decap_3 PHY_4670 ();
 sky130_fd_sc_hd__decap_3 PHY_4671 ();
 sky130_fd_sc_hd__decap_3 PHY_4672 ();
 sky130_fd_sc_hd__decap_3 PHY_4673 ();
 sky130_fd_sc_hd__decap_3 PHY_4674 ();
 sky130_fd_sc_hd__decap_3 PHY_4675 ();
 sky130_fd_sc_hd__decap_3 PHY_4676 ();
 sky130_fd_sc_hd__decap_3 PHY_4677 ();
 sky130_fd_sc_hd__decap_3 PHY_4678 ();
 sky130_fd_sc_hd__decap_3 PHY_4679 ();
 sky130_fd_sc_hd__decap_3 PHY_4680 ();
 sky130_fd_sc_hd__decap_3 PHY_4681 ();
 sky130_fd_sc_hd__decap_3 PHY_4682 ();
 sky130_fd_sc_hd__decap_3 PHY_4683 ();
 sky130_fd_sc_hd__decap_3 PHY_4684 ();
 sky130_fd_sc_hd__decap_3 PHY_4685 ();
 sky130_fd_sc_hd__decap_3 PHY_4686 ();
 sky130_fd_sc_hd__decap_3 PHY_4687 ();
 sky130_fd_sc_hd__decap_3 PHY_4688 ();
 sky130_fd_sc_hd__decap_3 PHY_4689 ();
 sky130_fd_sc_hd__decap_3 PHY_4690 ();
 sky130_fd_sc_hd__decap_3 PHY_4691 ();
 sky130_fd_sc_hd__decap_3 PHY_4692 ();
 sky130_fd_sc_hd__decap_3 PHY_4693 ();
 sky130_fd_sc_hd__decap_3 PHY_4694 ();
 sky130_fd_sc_hd__decap_3 PHY_4695 ();
 sky130_fd_sc_hd__decap_3 PHY_4696 ();
 sky130_fd_sc_hd__decap_3 PHY_4697 ();
 sky130_fd_sc_hd__decap_3 PHY_4698 ();
 sky130_fd_sc_hd__decap_3 PHY_4699 ();
 sky130_fd_sc_hd__decap_3 PHY_4700 ();
 sky130_fd_sc_hd__decap_3 PHY_4701 ();
 sky130_fd_sc_hd__decap_3 PHY_4702 ();
 sky130_fd_sc_hd__decap_3 PHY_4703 ();
 sky130_fd_sc_hd__decap_3 PHY_4704 ();
 sky130_fd_sc_hd__decap_3 PHY_4705 ();
 sky130_fd_sc_hd__decap_3 PHY_4706 ();
 sky130_fd_sc_hd__decap_3 PHY_4707 ();
 sky130_fd_sc_hd__decap_3 PHY_4708 ();
 sky130_fd_sc_hd__decap_3 PHY_4709 ();
 sky130_fd_sc_hd__decap_3 PHY_4710 ();
 sky130_fd_sc_hd__decap_3 PHY_4711 ();
 sky130_fd_sc_hd__decap_3 PHY_4712 ();
 sky130_fd_sc_hd__decap_3 PHY_4713 ();
 sky130_fd_sc_hd__decap_3 PHY_4714 ();
 sky130_fd_sc_hd__decap_3 PHY_4715 ();
 sky130_fd_sc_hd__decap_3 PHY_4716 ();
 sky130_fd_sc_hd__decap_3 PHY_4717 ();
 sky130_fd_sc_hd__decap_3 PHY_4718 ();
 sky130_fd_sc_hd__decap_3 PHY_4719 ();
 sky130_fd_sc_hd__decap_3 PHY_4720 ();
 sky130_fd_sc_hd__decap_3 PHY_4721 ();
 sky130_fd_sc_hd__decap_3 PHY_4722 ();
 sky130_fd_sc_hd__decap_3 PHY_4723 ();
 sky130_fd_sc_hd__decap_3 PHY_4724 ();
 sky130_fd_sc_hd__decap_3 PHY_4725 ();
 sky130_fd_sc_hd__decap_3 PHY_4726 ();
 sky130_fd_sc_hd__decap_3 PHY_4727 ();
 sky130_fd_sc_hd__decap_3 PHY_4728 ();
 sky130_fd_sc_hd__decap_3 PHY_4729 ();
 sky130_fd_sc_hd__decap_3 PHY_4730 ();
 sky130_fd_sc_hd__decap_3 PHY_4731 ();
 sky130_fd_sc_hd__decap_3 PHY_4732 ();
 sky130_fd_sc_hd__decap_3 PHY_4733 ();
 sky130_fd_sc_hd__decap_3 PHY_4734 ();
 sky130_fd_sc_hd__decap_3 PHY_4735 ();
 sky130_fd_sc_hd__decap_3 PHY_4736 ();
 sky130_fd_sc_hd__decap_3 PHY_4737 ();
 sky130_fd_sc_hd__decap_3 PHY_4738 ();
 sky130_fd_sc_hd__decap_3 PHY_4739 ();
 sky130_fd_sc_hd__decap_3 PHY_4740 ();
 sky130_fd_sc_hd__decap_3 PHY_4741 ();
 sky130_fd_sc_hd__decap_3 PHY_4742 ();
 sky130_fd_sc_hd__decap_3 PHY_4743 ();
 sky130_fd_sc_hd__decap_3 PHY_4744 ();
 sky130_fd_sc_hd__decap_3 PHY_4745 ();
 sky130_fd_sc_hd__decap_3 PHY_4746 ();
 sky130_fd_sc_hd__decap_3 PHY_4747 ();
 sky130_fd_sc_hd__decap_3 PHY_4748 ();
 sky130_fd_sc_hd__decap_3 PHY_4749 ();
 sky130_fd_sc_hd__decap_3 PHY_4750 ();
 sky130_fd_sc_hd__decap_3 PHY_4751 ();
 sky130_fd_sc_hd__decap_3 PHY_4752 ();
 sky130_fd_sc_hd__decap_3 PHY_4753 ();
 sky130_fd_sc_hd__decap_3 PHY_4754 ();
 sky130_fd_sc_hd__decap_3 PHY_4755 ();
 sky130_fd_sc_hd__decap_3 PHY_4756 ();
 sky130_fd_sc_hd__decap_3 PHY_4757 ();
 sky130_fd_sc_hd__decap_3 PHY_4758 ();
 sky130_fd_sc_hd__decap_3 PHY_4759 ();
 sky130_fd_sc_hd__decap_3 PHY_4760 ();
 sky130_fd_sc_hd__decap_3 PHY_4761 ();
 sky130_fd_sc_hd__decap_3 PHY_4762 ();
 sky130_fd_sc_hd__decap_3 PHY_4763 ();
 sky130_fd_sc_hd__decap_3 PHY_4764 ();
 sky130_fd_sc_hd__decap_3 PHY_4765 ();
 sky130_fd_sc_hd__decap_3 PHY_4766 ();
 sky130_fd_sc_hd__decap_3 PHY_4767 ();
 sky130_fd_sc_hd__decap_3 PHY_4768 ();
 sky130_fd_sc_hd__decap_3 PHY_4769 ();
 sky130_fd_sc_hd__decap_3 PHY_4770 ();
 sky130_fd_sc_hd__decap_3 PHY_4771 ();
 sky130_fd_sc_hd__decap_3 PHY_4772 ();
 sky130_fd_sc_hd__decap_3 PHY_4773 ();
 sky130_fd_sc_hd__decap_3 PHY_4774 ();
 sky130_fd_sc_hd__decap_3 PHY_4775 ();
 sky130_fd_sc_hd__decap_3 PHY_4776 ();
 sky130_fd_sc_hd__decap_3 PHY_4777 ();
 sky130_fd_sc_hd__decap_3 PHY_4778 ();
 sky130_fd_sc_hd__decap_3 PHY_4779 ();
 sky130_fd_sc_hd__decap_3 PHY_4780 ();
 sky130_fd_sc_hd__decap_3 PHY_4781 ();
 sky130_fd_sc_hd__decap_3 PHY_4782 ();
 sky130_fd_sc_hd__decap_3 PHY_4783 ();
 sky130_fd_sc_hd__decap_3 PHY_4784 ();
 sky130_fd_sc_hd__decap_3 PHY_4785 ();
 sky130_fd_sc_hd__decap_3 PHY_4786 ();
 sky130_fd_sc_hd__decap_3 PHY_4787 ();
 sky130_fd_sc_hd__decap_3 PHY_4788 ();
 sky130_fd_sc_hd__decap_3 PHY_4789 ();
 sky130_fd_sc_hd__decap_3 PHY_4790 ();
 sky130_fd_sc_hd__decap_3 PHY_4791 ();
 sky130_fd_sc_hd__decap_3 PHY_4792 ();
 sky130_fd_sc_hd__decap_3 PHY_4793 ();
 sky130_fd_sc_hd__decap_3 PHY_4794 ();
 sky130_fd_sc_hd__decap_3 PHY_4795 ();
 sky130_fd_sc_hd__decap_3 PHY_4796 ();
 sky130_fd_sc_hd__decap_3 PHY_4797 ();
 sky130_fd_sc_hd__decap_3 PHY_4798 ();
 sky130_fd_sc_hd__decap_3 PHY_4799 ();
 sky130_fd_sc_hd__decap_3 PHY_4800 ();
 sky130_fd_sc_hd__decap_3 PHY_4801 ();
 sky130_fd_sc_hd__decap_3 PHY_4802 ();
 sky130_fd_sc_hd__decap_3 PHY_4803 ();
 sky130_fd_sc_hd__decap_3 PHY_4804 ();
 sky130_fd_sc_hd__decap_3 PHY_4805 ();
 sky130_fd_sc_hd__decap_3 PHY_4806 ();
 sky130_fd_sc_hd__decap_3 PHY_4807 ();
 sky130_fd_sc_hd__decap_3 PHY_4808 ();
 sky130_fd_sc_hd__decap_3 PHY_4809 ();
 sky130_fd_sc_hd__decap_3 PHY_4810 ();
 sky130_fd_sc_hd__decap_3 PHY_4811 ();
 sky130_fd_sc_hd__decap_3 PHY_4812 ();
 sky130_fd_sc_hd__decap_3 PHY_4813 ();
 sky130_fd_sc_hd__decap_3 PHY_4814 ();
 sky130_fd_sc_hd__decap_3 PHY_4815 ();
 sky130_fd_sc_hd__decap_3 PHY_4816 ();
 sky130_fd_sc_hd__decap_3 PHY_4817 ();
 sky130_fd_sc_hd__decap_3 PHY_4818 ();
 sky130_fd_sc_hd__decap_3 PHY_4819 ();
 sky130_fd_sc_hd__decap_3 PHY_4820 ();
 sky130_fd_sc_hd__decap_3 PHY_4821 ();
 sky130_fd_sc_hd__decap_3 PHY_4822 ();
 sky130_fd_sc_hd__decap_3 PHY_4823 ();
 sky130_fd_sc_hd__decap_3 PHY_4824 ();
 sky130_fd_sc_hd__decap_3 PHY_4825 ();
 sky130_fd_sc_hd__decap_3 PHY_4826 ();
 sky130_fd_sc_hd__decap_3 PHY_4827 ();
 sky130_fd_sc_hd__decap_3 PHY_4828 ();
 sky130_fd_sc_hd__decap_3 PHY_4829 ();
 sky130_fd_sc_hd__decap_3 PHY_4830 ();
 sky130_fd_sc_hd__decap_3 PHY_4831 ();
 sky130_fd_sc_hd__decap_3 PHY_4832 ();
 sky130_fd_sc_hd__decap_3 PHY_4833 ();
 sky130_fd_sc_hd__decap_3 PHY_4834 ();
 sky130_fd_sc_hd__decap_3 PHY_4835 ();
 sky130_fd_sc_hd__decap_3 PHY_4836 ();
 sky130_fd_sc_hd__decap_3 PHY_4837 ();
 sky130_fd_sc_hd__decap_3 PHY_4838 ();
 sky130_fd_sc_hd__decap_3 PHY_4839 ();
 sky130_fd_sc_hd__decap_3 PHY_4840 ();
 sky130_fd_sc_hd__decap_3 PHY_4841 ();
 sky130_fd_sc_hd__decap_3 PHY_4842 ();
 sky130_fd_sc_hd__decap_3 PHY_4843 ();
 sky130_fd_sc_hd__decap_3 PHY_4844 ();
 sky130_fd_sc_hd__decap_3 PHY_4845 ();
 sky130_fd_sc_hd__decap_3 PHY_4846 ();
 sky130_fd_sc_hd__decap_3 PHY_4847 ();
 sky130_fd_sc_hd__decap_3 PHY_4848 ();
 sky130_fd_sc_hd__decap_3 PHY_4849 ();
 sky130_fd_sc_hd__decap_3 PHY_4850 ();
 sky130_fd_sc_hd__decap_3 PHY_4851 ();
 sky130_fd_sc_hd__decap_3 PHY_4852 ();
 sky130_fd_sc_hd__decap_3 PHY_4853 ();
 sky130_fd_sc_hd__decap_3 PHY_4854 ();
 sky130_fd_sc_hd__decap_3 PHY_4855 ();
 sky130_fd_sc_hd__decap_3 PHY_4856 ();
 sky130_fd_sc_hd__decap_3 PHY_4857 ();
 sky130_fd_sc_hd__decap_3 PHY_4858 ();
 sky130_fd_sc_hd__decap_3 PHY_4859 ();
 sky130_fd_sc_hd__decap_3 PHY_4860 ();
 sky130_fd_sc_hd__decap_3 PHY_4861 ();
 sky130_fd_sc_hd__decap_3 PHY_4862 ();
 sky130_fd_sc_hd__decap_3 PHY_4863 ();
 sky130_fd_sc_hd__decap_3 PHY_4864 ();
 sky130_fd_sc_hd__decap_3 PHY_4865 ();
 sky130_fd_sc_hd__decap_3 PHY_4866 ();
 sky130_fd_sc_hd__decap_3 PHY_4867 ();
 sky130_fd_sc_hd__decap_3 PHY_4868 ();
 sky130_fd_sc_hd__decap_3 PHY_4869 ();
 sky130_fd_sc_hd__decap_3 PHY_4870 ();
 sky130_fd_sc_hd__decap_3 PHY_4871 ();
 sky130_fd_sc_hd__decap_3 PHY_4872 ();
 sky130_fd_sc_hd__decap_3 PHY_4873 ();
 sky130_fd_sc_hd__decap_3 PHY_4874 ();
 sky130_fd_sc_hd__decap_3 PHY_4875 ();
 sky130_fd_sc_hd__decap_3 PHY_4876 ();
 sky130_fd_sc_hd__decap_3 PHY_4877 ();
 sky130_fd_sc_hd__decap_3 PHY_4878 ();
 sky130_fd_sc_hd__decap_3 PHY_4879 ();
 sky130_fd_sc_hd__decap_3 PHY_4880 ();
 sky130_fd_sc_hd__decap_3 PHY_4881 ();
 sky130_fd_sc_hd__decap_3 PHY_4882 ();
 sky130_fd_sc_hd__decap_3 PHY_4883 ();
 sky130_fd_sc_hd__decap_3 PHY_4884 ();
 sky130_fd_sc_hd__decap_3 PHY_4885 ();
 sky130_fd_sc_hd__decap_3 PHY_4886 ();
 sky130_fd_sc_hd__decap_3 PHY_4887 ();
 sky130_fd_sc_hd__decap_3 PHY_4888 ();
 sky130_fd_sc_hd__decap_3 PHY_4889 ();
 sky130_fd_sc_hd__decap_3 PHY_4890 ();
 sky130_fd_sc_hd__decap_3 PHY_4891 ();
 sky130_fd_sc_hd__decap_3 PHY_4892 ();
 sky130_fd_sc_hd__decap_3 PHY_4893 ();
 sky130_fd_sc_hd__decap_3 PHY_4894 ();
 sky130_fd_sc_hd__decap_3 PHY_4895 ();
 sky130_fd_sc_hd__decap_3 PHY_4896 ();
 sky130_fd_sc_hd__decap_3 PHY_4897 ();
 sky130_fd_sc_hd__decap_3 PHY_4898 ();
 sky130_fd_sc_hd__decap_3 PHY_4899 ();
 sky130_fd_sc_hd__decap_3 PHY_4900 ();
 sky130_fd_sc_hd__decap_3 PHY_4901 ();
 sky130_fd_sc_hd__decap_3 PHY_4902 ();
 sky130_fd_sc_hd__decap_3 PHY_4903 ();
 sky130_fd_sc_hd__decap_3 PHY_4904 ();
 sky130_fd_sc_hd__decap_3 PHY_4905 ();
 sky130_fd_sc_hd__decap_3 PHY_4906 ();
 sky130_fd_sc_hd__decap_3 PHY_4907 ();
 sky130_fd_sc_hd__decap_3 PHY_4908 ();
 sky130_fd_sc_hd__decap_3 PHY_4909 ();
 sky130_fd_sc_hd__decap_3 PHY_4910 ();
 sky130_fd_sc_hd__decap_3 PHY_4911 ();
 sky130_fd_sc_hd__decap_3 PHY_4912 ();
 sky130_fd_sc_hd__decap_3 PHY_4913 ();
 sky130_fd_sc_hd__decap_3 PHY_4914 ();
 sky130_fd_sc_hd__decap_3 PHY_4915 ();
 sky130_fd_sc_hd__decap_3 PHY_4916 ();
 sky130_fd_sc_hd__decap_3 PHY_4917 ();
 sky130_fd_sc_hd__decap_3 PHY_4918 ();
 sky130_fd_sc_hd__decap_3 PHY_4919 ();
 sky130_fd_sc_hd__decap_3 PHY_4920 ();
 sky130_fd_sc_hd__decap_3 PHY_4921 ();
 sky130_fd_sc_hd__decap_3 PHY_4922 ();
 sky130_fd_sc_hd__decap_3 PHY_4923 ();
 sky130_fd_sc_hd__decap_3 PHY_4924 ();
 sky130_fd_sc_hd__decap_3 PHY_4925 ();
 sky130_fd_sc_hd__decap_3 PHY_4926 ();
 sky130_fd_sc_hd__decap_3 PHY_4927 ();
 sky130_fd_sc_hd__decap_3 PHY_4928 ();
 sky130_fd_sc_hd__decap_3 PHY_4929 ();
 sky130_fd_sc_hd__decap_3 PHY_4930 ();
 sky130_fd_sc_hd__decap_3 PHY_4931 ();
 sky130_fd_sc_hd__decap_3 PHY_4932 ();
 sky130_fd_sc_hd__decap_3 PHY_4933 ();
 sky130_fd_sc_hd__decap_3 PHY_4934 ();
 sky130_fd_sc_hd__decap_3 PHY_4935 ();
 sky130_fd_sc_hd__decap_3 PHY_4936 ();
 sky130_fd_sc_hd__decap_3 PHY_4937 ();
 sky130_fd_sc_hd__decap_3 PHY_4938 ();
 sky130_fd_sc_hd__decap_3 PHY_4939 ();
 sky130_fd_sc_hd__decap_3 PHY_4940 ();
 sky130_fd_sc_hd__decap_3 PHY_4941 ();
 sky130_fd_sc_hd__decap_3 PHY_4942 ();
 sky130_fd_sc_hd__decap_3 PHY_4943 ();
 sky130_fd_sc_hd__decap_3 PHY_4944 ();
 sky130_fd_sc_hd__decap_3 PHY_4945 ();
 sky130_fd_sc_hd__decap_3 PHY_4946 ();
 sky130_fd_sc_hd__decap_3 PHY_4947 ();
 sky130_fd_sc_hd__decap_3 PHY_4948 ();
 sky130_fd_sc_hd__decap_3 PHY_4949 ();
 sky130_fd_sc_hd__decap_3 PHY_4950 ();
 sky130_fd_sc_hd__decap_3 PHY_4951 ();
 sky130_fd_sc_hd__decap_3 PHY_4952 ();
 sky130_fd_sc_hd__decap_3 PHY_4953 ();
 sky130_fd_sc_hd__decap_3 PHY_4954 ();
 sky130_fd_sc_hd__decap_3 PHY_4955 ();
 sky130_fd_sc_hd__decap_3 PHY_4956 ();
 sky130_fd_sc_hd__decap_3 PHY_4957 ();
 sky130_fd_sc_hd__decap_3 PHY_4958 ();
 sky130_fd_sc_hd__decap_3 PHY_4959 ();
 sky130_fd_sc_hd__decap_3 PHY_4960 ();
 sky130_fd_sc_hd__decap_3 PHY_4961 ();
 sky130_fd_sc_hd__decap_3 PHY_4962 ();
 sky130_fd_sc_hd__decap_3 PHY_4963 ();
 sky130_fd_sc_hd__decap_3 PHY_4964 ();
 sky130_fd_sc_hd__decap_3 PHY_4965 ();
 sky130_fd_sc_hd__decap_3 PHY_4966 ();
 sky130_fd_sc_hd__decap_3 PHY_4967 ();
 sky130_fd_sc_hd__decap_3 PHY_4968 ();
 sky130_fd_sc_hd__decap_3 PHY_4969 ();
 sky130_fd_sc_hd__decap_3 PHY_4970 ();
 sky130_fd_sc_hd__decap_3 PHY_4971 ();
 sky130_fd_sc_hd__decap_3 PHY_4972 ();
 sky130_fd_sc_hd__decap_3 PHY_4973 ();
 sky130_fd_sc_hd__decap_3 PHY_4974 ();
 sky130_fd_sc_hd__decap_3 PHY_4975 ();
 sky130_fd_sc_hd__decap_3 PHY_4976 ();
 sky130_fd_sc_hd__decap_3 PHY_4977 ();
 sky130_fd_sc_hd__decap_3 PHY_4978 ();
 sky130_fd_sc_hd__decap_3 PHY_4979 ();
 sky130_fd_sc_hd__decap_3 PHY_4980 ();
 sky130_fd_sc_hd__decap_3 PHY_4981 ();
 sky130_fd_sc_hd__decap_3 PHY_4982 ();
 sky130_fd_sc_hd__decap_3 PHY_4983 ();
 sky130_fd_sc_hd__decap_3 PHY_4984 ();
 sky130_fd_sc_hd__decap_3 PHY_4985 ();
 sky130_fd_sc_hd__decap_3 PHY_4986 ();
 sky130_fd_sc_hd__decap_3 PHY_4987 ();
 sky130_fd_sc_hd__decap_3 PHY_4988 ();
 sky130_fd_sc_hd__decap_3 PHY_4989 ();
 sky130_fd_sc_hd__decap_3 PHY_4990 ();
 sky130_fd_sc_hd__decap_3 PHY_4991 ();
 sky130_fd_sc_hd__decap_3 PHY_4992 ();
 sky130_fd_sc_hd__decap_3 PHY_4993 ();
 sky130_fd_sc_hd__decap_3 PHY_4994 ();
 sky130_fd_sc_hd__decap_3 PHY_4995 ();
 sky130_fd_sc_hd__decap_3 PHY_4996 ();
 sky130_fd_sc_hd__decap_3 PHY_4997 ();
 sky130_fd_sc_hd__decap_3 PHY_4998 ();
 sky130_fd_sc_hd__decap_3 PHY_4999 ();
 sky130_fd_sc_hd__decap_3 PHY_5000 ();
 sky130_fd_sc_hd__decap_3 PHY_5001 ();
 sky130_fd_sc_hd__decap_3 PHY_5002 ();
 sky130_fd_sc_hd__decap_3 PHY_5003 ();
 sky130_fd_sc_hd__decap_3 PHY_5004 ();
 sky130_fd_sc_hd__decap_3 PHY_5005 ();
 sky130_fd_sc_hd__decap_3 PHY_5006 ();
 sky130_fd_sc_hd__decap_3 PHY_5007 ();
 sky130_fd_sc_hd__decap_3 PHY_5008 ();
 sky130_fd_sc_hd__decap_3 PHY_5009 ();
 sky130_fd_sc_hd__decap_3 PHY_5010 ();
 sky130_fd_sc_hd__decap_3 PHY_5011 ();
 sky130_fd_sc_hd__decap_3 PHY_5012 ();
 sky130_fd_sc_hd__decap_3 PHY_5013 ();
 sky130_fd_sc_hd__decap_3 PHY_5014 ();
 sky130_fd_sc_hd__decap_3 PHY_5015 ();
 sky130_fd_sc_hd__decap_3 PHY_5016 ();
 sky130_fd_sc_hd__decap_3 PHY_5017 ();
 sky130_fd_sc_hd__decap_3 PHY_5018 ();
 sky130_fd_sc_hd__decap_3 PHY_5019 ();
 sky130_fd_sc_hd__decap_3 PHY_5020 ();
 sky130_fd_sc_hd__decap_3 PHY_5021 ();
 sky130_fd_sc_hd__decap_3 PHY_5022 ();
 sky130_fd_sc_hd__decap_3 PHY_5023 ();
 sky130_fd_sc_hd__decap_3 PHY_5024 ();
 sky130_fd_sc_hd__decap_3 PHY_5025 ();
 sky130_fd_sc_hd__decap_3 PHY_5026 ();
 sky130_fd_sc_hd__decap_3 PHY_5027 ();
 sky130_fd_sc_hd__decap_3 PHY_5028 ();
 sky130_fd_sc_hd__decap_3 PHY_5029 ();
 sky130_fd_sc_hd__decap_3 PHY_5030 ();
 sky130_fd_sc_hd__decap_3 PHY_5031 ();
 sky130_fd_sc_hd__decap_3 PHY_5032 ();
 sky130_fd_sc_hd__decap_3 PHY_5033 ();
 sky130_fd_sc_hd__decap_3 PHY_5034 ();
 sky130_fd_sc_hd__decap_3 PHY_5035 ();
 sky130_fd_sc_hd__decap_3 PHY_5036 ();
 sky130_fd_sc_hd__decap_3 PHY_5037 ();
 sky130_fd_sc_hd__decap_3 PHY_5038 ();
 sky130_fd_sc_hd__decap_3 PHY_5039 ();
 sky130_fd_sc_hd__decap_3 PHY_5040 ();
 sky130_fd_sc_hd__decap_3 PHY_5041 ();
 sky130_fd_sc_hd__decap_3 PHY_5042 ();
 sky130_fd_sc_hd__decap_3 PHY_5043 ();
 sky130_fd_sc_hd__decap_3 PHY_5044 ();
 sky130_fd_sc_hd__decap_3 PHY_5045 ();
 sky130_fd_sc_hd__decap_3 PHY_5046 ();
 sky130_fd_sc_hd__decap_3 PHY_5047 ();
 sky130_fd_sc_hd__decap_3 PHY_5048 ();
 sky130_fd_sc_hd__decap_3 PHY_5049 ();
 sky130_fd_sc_hd__decap_3 PHY_5050 ();
 sky130_fd_sc_hd__decap_3 PHY_5051 ();
 sky130_fd_sc_hd__decap_3 PHY_5052 ();
 sky130_fd_sc_hd__decap_3 PHY_5053 ();
 sky130_fd_sc_hd__decap_3 PHY_5054 ();
 sky130_fd_sc_hd__decap_3 PHY_5055 ();
 sky130_fd_sc_hd__decap_3 PHY_5056 ();
 sky130_fd_sc_hd__decap_3 PHY_5057 ();
 sky130_fd_sc_hd__decap_3 PHY_5058 ();
 sky130_fd_sc_hd__decap_3 PHY_5059 ();
 sky130_fd_sc_hd__decap_3 PHY_5060 ();
 sky130_fd_sc_hd__decap_3 PHY_5061 ();
 sky130_fd_sc_hd__decap_3 PHY_5062 ();
 sky130_fd_sc_hd__decap_3 PHY_5063 ();
 sky130_fd_sc_hd__decap_3 PHY_5064 ();
 sky130_fd_sc_hd__decap_3 PHY_5065 ();
 sky130_fd_sc_hd__decap_3 PHY_5066 ();
 sky130_fd_sc_hd__decap_3 PHY_5067 ();
 sky130_fd_sc_hd__decap_3 PHY_5068 ();
 sky130_fd_sc_hd__decap_3 PHY_5069 ();
 sky130_fd_sc_hd__decap_3 PHY_5070 ();
 sky130_fd_sc_hd__decap_3 PHY_5071 ();
 sky130_fd_sc_hd__decap_3 PHY_5072 ();
 sky130_fd_sc_hd__decap_3 PHY_5073 ();
 sky130_fd_sc_hd__decap_3 PHY_5074 ();
 sky130_fd_sc_hd__decap_3 PHY_5075 ();
 sky130_fd_sc_hd__decap_3 PHY_5076 ();
 sky130_fd_sc_hd__decap_3 PHY_5077 ();
 sky130_fd_sc_hd__decap_3 PHY_5078 ();
 sky130_fd_sc_hd__decap_3 PHY_5079 ();
 sky130_fd_sc_hd__decap_3 PHY_5080 ();
 sky130_fd_sc_hd__decap_3 PHY_5081 ();
 sky130_fd_sc_hd__decap_3 PHY_5082 ();
 sky130_fd_sc_hd__decap_3 PHY_5083 ();
 sky130_fd_sc_hd__decap_3 PHY_5084 ();
 sky130_fd_sc_hd__decap_3 PHY_5085 ();
 sky130_fd_sc_hd__decap_3 PHY_5086 ();
 sky130_fd_sc_hd__decap_3 PHY_5087 ();
 sky130_fd_sc_hd__decap_3 PHY_5088 ();
 sky130_fd_sc_hd__decap_3 PHY_5089 ();
 sky130_fd_sc_hd__decap_3 PHY_5090 ();
 sky130_fd_sc_hd__decap_3 PHY_5091 ();
 sky130_fd_sc_hd__decap_3 PHY_5092 ();
 sky130_fd_sc_hd__decap_3 PHY_5093 ();
 sky130_fd_sc_hd__decap_3 PHY_5094 ();
 sky130_fd_sc_hd__decap_3 PHY_5095 ();
 sky130_fd_sc_hd__decap_3 PHY_5096 ();
 sky130_fd_sc_hd__decap_3 PHY_5097 ();
 sky130_fd_sc_hd__decap_3 PHY_5098 ();
 sky130_fd_sc_hd__decap_3 PHY_5099 ();
 sky130_fd_sc_hd__decap_3 PHY_5100 ();
 sky130_fd_sc_hd__decap_3 PHY_5101 ();
 sky130_fd_sc_hd__decap_3 PHY_5102 ();
 sky130_fd_sc_hd__decap_3 PHY_5103 ();
 sky130_fd_sc_hd__decap_3 PHY_5104 ();
 sky130_fd_sc_hd__decap_3 PHY_5105 ();
 sky130_fd_sc_hd__decap_3 PHY_5106 ();
 sky130_fd_sc_hd__decap_3 PHY_5107 ();
 sky130_fd_sc_hd__decap_3 PHY_5108 ();
 sky130_fd_sc_hd__decap_3 PHY_5109 ();
 sky130_fd_sc_hd__decap_3 PHY_5110 ();
 sky130_fd_sc_hd__decap_3 PHY_5111 ();
 sky130_fd_sc_hd__decap_3 PHY_5112 ();
 sky130_fd_sc_hd__decap_3 PHY_5113 ();
 sky130_fd_sc_hd__decap_3 PHY_5114 ();
 sky130_fd_sc_hd__decap_3 PHY_5115 ();
 sky130_fd_sc_hd__decap_3 PHY_5116 ();
 sky130_fd_sc_hd__decap_3 PHY_5117 ();
 sky130_fd_sc_hd__decap_3 PHY_5118 ();
 sky130_fd_sc_hd__decap_3 PHY_5119 ();
 sky130_fd_sc_hd__decap_3 PHY_5120 ();
 sky130_fd_sc_hd__decap_3 PHY_5121 ();
 sky130_fd_sc_hd__decap_3 PHY_5122 ();
 sky130_fd_sc_hd__decap_3 PHY_5123 ();
 sky130_fd_sc_hd__decap_3 PHY_5124 ();
 sky130_fd_sc_hd__decap_3 PHY_5125 ();
 sky130_fd_sc_hd__decap_3 PHY_5126 ();
 sky130_fd_sc_hd__decap_3 PHY_5127 ();
 sky130_fd_sc_hd__decap_3 PHY_5128 ();
 sky130_fd_sc_hd__decap_3 PHY_5129 ();
 sky130_fd_sc_hd__decap_3 PHY_5130 ();
 sky130_fd_sc_hd__decap_3 PHY_5131 ();
 sky130_fd_sc_hd__decap_3 PHY_5132 ();
 sky130_fd_sc_hd__decap_3 PHY_5133 ();
 sky130_fd_sc_hd__decap_3 PHY_5134 ();
 sky130_fd_sc_hd__decap_3 PHY_5135 ();
 sky130_fd_sc_hd__decap_3 PHY_5136 ();
 sky130_fd_sc_hd__decap_3 PHY_5137 ();
 sky130_fd_sc_hd__decap_3 PHY_5138 ();
 sky130_fd_sc_hd__decap_3 PHY_5139 ();
 sky130_fd_sc_hd__decap_3 PHY_5140 ();
 sky130_fd_sc_hd__decap_3 PHY_5141 ();
 sky130_fd_sc_hd__decap_3 PHY_5142 ();
 sky130_fd_sc_hd__decap_3 PHY_5143 ();
 sky130_fd_sc_hd__decap_3 PHY_5144 ();
 sky130_fd_sc_hd__decap_3 PHY_5145 ();
 sky130_fd_sc_hd__decap_3 PHY_5146 ();
 sky130_fd_sc_hd__decap_3 PHY_5147 ();
 sky130_fd_sc_hd__decap_3 PHY_5148 ();
 sky130_fd_sc_hd__decap_3 PHY_5149 ();
 sky130_fd_sc_hd__decap_3 PHY_5150 ();
 sky130_fd_sc_hd__decap_3 PHY_5151 ();
 sky130_fd_sc_hd__decap_3 PHY_5152 ();
 sky130_fd_sc_hd__decap_3 PHY_5153 ();
 sky130_fd_sc_hd__decap_3 PHY_5154 ();
 sky130_fd_sc_hd__decap_3 PHY_5155 ();
 sky130_fd_sc_hd__decap_3 PHY_5156 ();
 sky130_fd_sc_hd__decap_3 PHY_5157 ();
 sky130_fd_sc_hd__decap_3 PHY_5158 ();
 sky130_fd_sc_hd__decap_3 PHY_5159 ();
 sky130_fd_sc_hd__decap_3 PHY_5160 ();
 sky130_fd_sc_hd__decap_3 PHY_5161 ();
 sky130_fd_sc_hd__decap_3 PHY_5162 ();
 sky130_fd_sc_hd__decap_3 PHY_5163 ();
 sky130_fd_sc_hd__decap_3 PHY_5164 ();
 sky130_fd_sc_hd__decap_3 PHY_5165 ();
 sky130_fd_sc_hd__decap_3 PHY_5166 ();
 sky130_fd_sc_hd__decap_3 PHY_5167 ();
 sky130_fd_sc_hd__decap_3 PHY_5168 ();
 sky130_fd_sc_hd__decap_3 PHY_5169 ();
 sky130_fd_sc_hd__decap_3 PHY_5170 ();
 sky130_fd_sc_hd__decap_3 PHY_5171 ();
 sky130_fd_sc_hd__decap_3 PHY_5172 ();
 sky130_fd_sc_hd__decap_3 PHY_5173 ();
 sky130_fd_sc_hd__decap_3 PHY_5174 ();
 sky130_fd_sc_hd__decap_3 PHY_5175 ();
 sky130_fd_sc_hd__decap_3 PHY_5176 ();
 sky130_fd_sc_hd__decap_3 PHY_5177 ();
 sky130_fd_sc_hd__decap_3 PHY_5178 ();
 sky130_fd_sc_hd__decap_3 PHY_5179 ();
 sky130_fd_sc_hd__decap_3 PHY_5180 ();
 sky130_fd_sc_hd__decap_3 PHY_5181 ();
 sky130_fd_sc_hd__decap_3 PHY_5182 ();
 sky130_fd_sc_hd__decap_3 PHY_5183 ();
 sky130_fd_sc_hd__decap_3 PHY_5184 ();
 sky130_fd_sc_hd__decap_3 PHY_5185 ();
 sky130_fd_sc_hd__decap_3 PHY_5186 ();
 sky130_fd_sc_hd__decap_3 PHY_5187 ();
 sky130_fd_sc_hd__decap_3 PHY_5188 ();
 sky130_fd_sc_hd__decap_3 PHY_5189 ();
 sky130_fd_sc_hd__decap_3 PHY_5190 ();
 sky130_fd_sc_hd__decap_3 PHY_5191 ();
 sky130_fd_sc_hd__decap_3 PHY_5192 ();
 sky130_fd_sc_hd__decap_3 PHY_5193 ();
 sky130_fd_sc_hd__decap_3 PHY_5194 ();
 sky130_fd_sc_hd__decap_3 PHY_5195 ();
 sky130_fd_sc_hd__decap_3 PHY_5196 ();
 sky130_fd_sc_hd__decap_3 PHY_5197 ();
 sky130_fd_sc_hd__decap_3 PHY_5198 ();
 sky130_fd_sc_hd__decap_3 PHY_5199 ();
 sky130_fd_sc_hd__decap_3 PHY_5200 ();
 sky130_fd_sc_hd__decap_3 PHY_5201 ();
 sky130_fd_sc_hd__decap_3 PHY_5202 ();
 sky130_fd_sc_hd__decap_3 PHY_5203 ();
 sky130_fd_sc_hd__decap_3 PHY_5204 ();
 sky130_fd_sc_hd__decap_3 PHY_5205 ();
 sky130_fd_sc_hd__decap_3 PHY_5206 ();
 sky130_fd_sc_hd__decap_3 PHY_5207 ();
 sky130_fd_sc_hd__decap_3 PHY_5208 ();
 sky130_fd_sc_hd__decap_3 PHY_5209 ();
 sky130_fd_sc_hd__decap_3 PHY_5210 ();
 sky130_fd_sc_hd__decap_3 PHY_5211 ();
 sky130_fd_sc_hd__decap_3 PHY_5212 ();
 sky130_fd_sc_hd__decap_3 PHY_5213 ();
 sky130_fd_sc_hd__decap_3 PHY_5214 ();
 sky130_fd_sc_hd__decap_3 PHY_5215 ();
 sky130_fd_sc_hd__decap_3 PHY_5216 ();
 sky130_fd_sc_hd__decap_3 PHY_5217 ();
 sky130_fd_sc_hd__decap_3 PHY_5218 ();
 sky130_fd_sc_hd__decap_3 PHY_5219 ();
 sky130_fd_sc_hd__decap_3 PHY_5220 ();
 sky130_fd_sc_hd__decap_3 PHY_5221 ();
 sky130_fd_sc_hd__decap_3 PHY_5222 ();
 sky130_fd_sc_hd__decap_3 PHY_5223 ();
 sky130_fd_sc_hd__decap_3 PHY_5224 ();
 sky130_fd_sc_hd__decap_3 PHY_5225 ();
 sky130_fd_sc_hd__decap_3 PHY_5226 ();
 sky130_fd_sc_hd__decap_3 PHY_5227 ();
 sky130_fd_sc_hd__decap_3 PHY_5228 ();
 sky130_fd_sc_hd__decap_3 PHY_5229 ();
 sky130_fd_sc_hd__decap_3 PHY_5230 ();
 sky130_fd_sc_hd__decap_3 PHY_5231 ();
 sky130_fd_sc_hd__decap_3 PHY_5232 ();
 sky130_fd_sc_hd__decap_3 PHY_5233 ();
 sky130_fd_sc_hd__decap_3 PHY_5234 ();
 sky130_fd_sc_hd__decap_3 PHY_5235 ();
 sky130_fd_sc_hd__decap_3 PHY_5236 ();
 sky130_fd_sc_hd__decap_3 PHY_5237 ();
 sky130_fd_sc_hd__decap_3 PHY_5238 ();
 sky130_fd_sc_hd__decap_3 PHY_5239 ();
 sky130_fd_sc_hd__decap_3 PHY_5240 ();
 sky130_fd_sc_hd__decap_3 PHY_5241 ();
 sky130_fd_sc_hd__decap_3 PHY_5242 ();
 sky130_fd_sc_hd__decap_3 PHY_5243 ();
 sky130_fd_sc_hd__decap_3 PHY_5244 ();
 sky130_fd_sc_hd__decap_3 PHY_5245 ();
 sky130_fd_sc_hd__decap_3 PHY_5246 ();
 sky130_fd_sc_hd__decap_3 PHY_5247 ();
 sky130_fd_sc_hd__decap_3 PHY_5248 ();
 sky130_fd_sc_hd__decap_3 PHY_5249 ();
 sky130_fd_sc_hd__decap_3 PHY_5250 ();
 sky130_fd_sc_hd__decap_3 PHY_5251 ();
 sky130_fd_sc_hd__decap_3 PHY_5252 ();
 sky130_fd_sc_hd__decap_3 PHY_5253 ();
 sky130_fd_sc_hd__decap_3 PHY_5254 ();
 sky130_fd_sc_hd__decap_3 PHY_5255 ();
 sky130_fd_sc_hd__decap_3 PHY_5256 ();
 sky130_fd_sc_hd__decap_3 PHY_5257 ();
 sky130_fd_sc_hd__decap_3 PHY_5258 ();
 sky130_fd_sc_hd__decap_3 PHY_5259 ();
 sky130_fd_sc_hd__decap_3 PHY_5260 ();
 sky130_fd_sc_hd__decap_3 PHY_5261 ();
 sky130_fd_sc_hd__decap_3 PHY_5262 ();
 sky130_fd_sc_hd__decap_3 PHY_5263 ();
 sky130_fd_sc_hd__decap_3 PHY_5264 ();
 sky130_fd_sc_hd__decap_3 PHY_5265 ();
 sky130_fd_sc_hd__decap_3 PHY_5266 ();
 sky130_fd_sc_hd__decap_3 PHY_5267 ();
 sky130_fd_sc_hd__decap_3 PHY_5268 ();
 sky130_fd_sc_hd__decap_3 PHY_5269 ();
 sky130_fd_sc_hd__decap_3 PHY_5270 ();
 sky130_fd_sc_hd__decap_3 PHY_5271 ();
 sky130_fd_sc_hd__decap_3 PHY_5272 ();
 sky130_fd_sc_hd__decap_3 PHY_5273 ();
 sky130_fd_sc_hd__decap_3 PHY_5274 ();
 sky130_fd_sc_hd__decap_3 PHY_5275 ();
 sky130_fd_sc_hd__decap_3 PHY_5276 ();
 sky130_fd_sc_hd__decap_3 PHY_5277 ();
 sky130_fd_sc_hd__decap_3 PHY_5278 ();
 sky130_fd_sc_hd__decap_3 PHY_5279 ();
 sky130_fd_sc_hd__decap_3 PHY_5280 ();
 sky130_fd_sc_hd__decap_3 PHY_5281 ();
 sky130_fd_sc_hd__decap_3 PHY_5282 ();
 sky130_fd_sc_hd__decap_3 PHY_5283 ();
 sky130_fd_sc_hd__decap_3 PHY_5284 ();
 sky130_fd_sc_hd__decap_3 PHY_5285 ();
 sky130_fd_sc_hd__decap_3 PHY_5286 ();
 sky130_fd_sc_hd__decap_3 PHY_5287 ();
 sky130_fd_sc_hd__decap_3 PHY_5288 ();
 sky130_fd_sc_hd__decap_3 PHY_5289 ();
 sky130_fd_sc_hd__decap_3 PHY_5290 ();
 sky130_fd_sc_hd__decap_3 PHY_5291 ();
 sky130_fd_sc_hd__decap_3 PHY_5292 ();
 sky130_fd_sc_hd__decap_3 PHY_5293 ();
 sky130_fd_sc_hd__decap_3 PHY_5294 ();
 sky130_fd_sc_hd__decap_3 PHY_5295 ();
 sky130_fd_sc_hd__decap_3 PHY_5296 ();
 sky130_fd_sc_hd__decap_3 PHY_5297 ();
 sky130_fd_sc_hd__decap_3 PHY_5298 ();
 sky130_fd_sc_hd__decap_3 PHY_5299 ();
 sky130_fd_sc_hd__decap_3 PHY_5300 ();
 sky130_fd_sc_hd__decap_3 PHY_5301 ();
 sky130_fd_sc_hd__decap_3 PHY_5302 ();
 sky130_fd_sc_hd__decap_3 PHY_5303 ();
 sky130_fd_sc_hd__decap_3 PHY_5304 ();
 sky130_fd_sc_hd__decap_3 PHY_5305 ();
 sky130_fd_sc_hd__decap_3 PHY_5306 ();
 sky130_fd_sc_hd__decap_3 PHY_5307 ();
 sky130_fd_sc_hd__decap_3 PHY_5308 ();
 sky130_fd_sc_hd__decap_3 PHY_5309 ();
 sky130_fd_sc_hd__decap_3 PHY_5310 ();
 sky130_fd_sc_hd__decap_3 PHY_5311 ();
 sky130_fd_sc_hd__decap_3 PHY_5312 ();
 sky130_fd_sc_hd__decap_3 PHY_5313 ();
 sky130_fd_sc_hd__decap_3 PHY_5314 ();
 sky130_fd_sc_hd__decap_3 PHY_5315 ();
 sky130_fd_sc_hd__decap_3 PHY_5316 ();
 sky130_fd_sc_hd__decap_3 PHY_5317 ();
 sky130_fd_sc_hd__decap_3 PHY_5318 ();
 sky130_fd_sc_hd__decap_3 PHY_5319 ();
 sky130_fd_sc_hd__decap_3 PHY_5320 ();
 sky130_fd_sc_hd__decap_3 PHY_5321 ();
 sky130_fd_sc_hd__decap_3 PHY_5322 ();
 sky130_fd_sc_hd__decap_3 PHY_5323 ();
 sky130_fd_sc_hd__decap_3 PHY_5324 ();
 sky130_fd_sc_hd__decap_3 PHY_5325 ();
 sky130_fd_sc_hd__decap_3 PHY_5326 ();
 sky130_fd_sc_hd__decap_3 PHY_5327 ();
 sky130_fd_sc_hd__decap_3 PHY_5328 ();
 sky130_fd_sc_hd__decap_3 PHY_5329 ();
 sky130_fd_sc_hd__decap_3 PHY_5330 ();
 sky130_fd_sc_hd__decap_3 PHY_5331 ();
 sky130_fd_sc_hd__decap_3 PHY_5332 ();
 sky130_fd_sc_hd__decap_3 PHY_5333 ();
 sky130_fd_sc_hd__decap_3 PHY_5334 ();
 sky130_fd_sc_hd__decap_3 PHY_5335 ();
 sky130_fd_sc_hd__decap_3 PHY_5336 ();
 sky130_fd_sc_hd__decap_3 PHY_5337 ();
 sky130_fd_sc_hd__decap_3 PHY_5338 ();
 sky130_fd_sc_hd__decap_3 PHY_5339 ();
 sky130_fd_sc_hd__decap_3 PHY_5340 ();
 sky130_fd_sc_hd__decap_3 PHY_5341 ();
 sky130_fd_sc_hd__decap_3 PHY_5342 ();
 sky130_fd_sc_hd__decap_3 PHY_5343 ();
 sky130_fd_sc_hd__decap_3 PHY_5344 ();
 sky130_fd_sc_hd__decap_3 PHY_5345 ();
 sky130_fd_sc_hd__decap_3 PHY_5346 ();
 sky130_fd_sc_hd__decap_3 PHY_5347 ();
 sky130_fd_sc_hd__decap_3 PHY_5348 ();
 sky130_fd_sc_hd__decap_3 PHY_5349 ();
 sky130_fd_sc_hd__decap_3 PHY_5350 ();
 sky130_fd_sc_hd__decap_3 PHY_5351 ();
 sky130_fd_sc_hd__decap_3 PHY_5352 ();
 sky130_fd_sc_hd__decap_3 PHY_5353 ();
 sky130_fd_sc_hd__decap_3 PHY_5354 ();
 sky130_fd_sc_hd__decap_3 PHY_5355 ();
 sky130_fd_sc_hd__decap_3 PHY_5356 ();
 sky130_fd_sc_hd__decap_3 PHY_5357 ();
 sky130_fd_sc_hd__decap_3 PHY_5358 ();
 sky130_fd_sc_hd__decap_3 PHY_5359 ();
 sky130_fd_sc_hd__decap_3 PHY_5360 ();
 sky130_fd_sc_hd__decap_3 PHY_5361 ();
 sky130_fd_sc_hd__decap_3 PHY_5362 ();
 sky130_fd_sc_hd__decap_3 PHY_5363 ();
 sky130_fd_sc_hd__decap_3 PHY_5364 ();
 sky130_fd_sc_hd__decap_3 PHY_5365 ();
 sky130_fd_sc_hd__decap_3 PHY_5366 ();
 sky130_fd_sc_hd__decap_3 PHY_5367 ();
 sky130_fd_sc_hd__decap_3 PHY_5368 ();
 sky130_fd_sc_hd__decap_3 PHY_5369 ();
 sky130_fd_sc_hd__decap_3 PHY_5370 ();
 sky130_fd_sc_hd__decap_3 PHY_5371 ();
 sky130_fd_sc_hd__decap_3 PHY_5372 ();
 sky130_fd_sc_hd__decap_3 PHY_5373 ();
 sky130_fd_sc_hd__decap_3 PHY_5374 ();
 sky130_fd_sc_hd__decap_3 PHY_5375 ();
 sky130_fd_sc_hd__decap_3 PHY_5376 ();
 sky130_fd_sc_hd__decap_3 PHY_5377 ();
 sky130_fd_sc_hd__decap_3 PHY_5378 ();
 sky130_fd_sc_hd__decap_3 PHY_5379 ();
 sky130_fd_sc_hd__decap_3 PHY_5380 ();
 sky130_fd_sc_hd__decap_3 PHY_5381 ();
 sky130_fd_sc_hd__decap_3 PHY_5382 ();
 sky130_fd_sc_hd__decap_3 PHY_5383 ();
 sky130_fd_sc_hd__decap_3 PHY_5384 ();
 sky130_fd_sc_hd__decap_3 PHY_5385 ();
 sky130_fd_sc_hd__decap_3 PHY_5386 ();
 sky130_fd_sc_hd__decap_3 PHY_5387 ();
 sky130_fd_sc_hd__decap_3 PHY_5388 ();
 sky130_fd_sc_hd__decap_3 PHY_5389 ();
 sky130_fd_sc_hd__decap_3 PHY_5390 ();
 sky130_fd_sc_hd__decap_3 PHY_5391 ();
 sky130_fd_sc_hd__decap_3 PHY_5392 ();
 sky130_fd_sc_hd__decap_3 PHY_5393 ();
 sky130_fd_sc_hd__decap_3 PHY_5394 ();
 sky130_fd_sc_hd__decap_3 PHY_5395 ();
 sky130_fd_sc_hd__decap_3 PHY_5396 ();
 sky130_fd_sc_hd__decap_3 PHY_5397 ();
 sky130_fd_sc_hd__decap_3 PHY_5398 ();
 sky130_fd_sc_hd__decap_3 PHY_5399 ();
 sky130_fd_sc_hd__decap_3 PHY_5400 ();
 sky130_fd_sc_hd__decap_3 PHY_5401 ();
 sky130_fd_sc_hd__decap_3 PHY_5402 ();
 sky130_fd_sc_hd__decap_3 PHY_5403 ();
 sky130_fd_sc_hd__decap_3 PHY_5404 ();
 sky130_fd_sc_hd__decap_3 PHY_5405 ();
 sky130_fd_sc_hd__decap_3 PHY_5406 ();
 sky130_fd_sc_hd__decap_3 PHY_5407 ();
 sky130_fd_sc_hd__decap_3 PHY_5408 ();
 sky130_fd_sc_hd__decap_3 PHY_5409 ();
 sky130_fd_sc_hd__decap_3 PHY_5410 ();
 sky130_fd_sc_hd__decap_3 PHY_5411 ();
 sky130_fd_sc_hd__decap_3 PHY_5412 ();
 sky130_fd_sc_hd__decap_3 PHY_5413 ();
 sky130_fd_sc_hd__decap_3 PHY_5414 ();
 sky130_fd_sc_hd__decap_3 PHY_5415 ();
 sky130_fd_sc_hd__decap_3 PHY_5416 ();
 sky130_fd_sc_hd__decap_3 PHY_5417 ();
 sky130_fd_sc_hd__decap_3 PHY_5418 ();
 sky130_fd_sc_hd__decap_3 PHY_5419 ();
 sky130_fd_sc_hd__decap_3 PHY_5420 ();
 sky130_fd_sc_hd__decap_3 PHY_5421 ();
 sky130_fd_sc_hd__decap_3 PHY_5422 ();
 sky130_fd_sc_hd__decap_3 PHY_5423 ();
 sky130_fd_sc_hd__decap_3 PHY_5424 ();
 sky130_fd_sc_hd__decap_3 PHY_5425 ();
 sky130_fd_sc_hd__decap_3 PHY_5426 ();
 sky130_fd_sc_hd__decap_3 PHY_5427 ();
 sky130_fd_sc_hd__decap_3 PHY_5428 ();
 sky130_fd_sc_hd__decap_3 PHY_5429 ();
 sky130_fd_sc_hd__decap_3 PHY_5430 ();
 sky130_fd_sc_hd__decap_3 PHY_5431 ();
 sky130_fd_sc_hd__decap_3 PHY_5432 ();
 sky130_fd_sc_hd__decap_3 PHY_5433 ();
 sky130_fd_sc_hd__decap_3 PHY_5434 ();
 sky130_fd_sc_hd__decap_3 PHY_5435 ();
 sky130_fd_sc_hd__decap_3 PHY_5436 ();
 sky130_fd_sc_hd__decap_3 PHY_5437 ();
 sky130_fd_sc_hd__decap_3 PHY_5438 ();
 sky130_fd_sc_hd__decap_3 PHY_5439 ();
 sky130_fd_sc_hd__decap_3 PHY_5440 ();
 sky130_fd_sc_hd__decap_3 PHY_5441 ();
 sky130_fd_sc_hd__decap_3 PHY_5442 ();
 sky130_fd_sc_hd__decap_3 PHY_5443 ();
 sky130_fd_sc_hd__decap_3 PHY_5444 ();
 sky130_fd_sc_hd__decap_3 PHY_5445 ();
 sky130_fd_sc_hd__decap_3 PHY_5446 ();
 sky130_fd_sc_hd__decap_3 PHY_5447 ();
 sky130_fd_sc_hd__decap_3 PHY_5448 ();
 sky130_fd_sc_hd__decap_3 PHY_5449 ();
 sky130_fd_sc_hd__decap_3 PHY_5450 ();
 sky130_fd_sc_hd__decap_3 PHY_5451 ();
 sky130_fd_sc_hd__decap_3 PHY_5452 ();
 sky130_fd_sc_hd__decap_3 PHY_5453 ();
 sky130_fd_sc_hd__decap_3 PHY_5454 ();
 sky130_fd_sc_hd__decap_3 PHY_5455 ();
 sky130_fd_sc_hd__decap_3 PHY_5456 ();
 sky130_fd_sc_hd__decap_3 PHY_5457 ();
 sky130_fd_sc_hd__decap_3 PHY_5458 ();
 sky130_fd_sc_hd__decap_3 PHY_5459 ();
 sky130_fd_sc_hd__decap_3 PHY_5460 ();
 sky130_fd_sc_hd__decap_3 PHY_5461 ();
 sky130_fd_sc_hd__decap_3 PHY_5462 ();
 sky130_fd_sc_hd__decap_3 PHY_5463 ();
 sky130_fd_sc_hd__decap_3 PHY_5464 ();
 sky130_fd_sc_hd__decap_3 PHY_5465 ();
 sky130_fd_sc_hd__decap_3 PHY_5466 ();
 sky130_fd_sc_hd__decap_3 PHY_5467 ();
 sky130_fd_sc_hd__decap_3 PHY_5468 ();
 sky130_fd_sc_hd__decap_3 PHY_5469 ();
 sky130_fd_sc_hd__decap_3 PHY_5470 ();
 sky130_fd_sc_hd__decap_3 PHY_5471 ();
 sky130_fd_sc_hd__decap_3 PHY_5472 ();
 sky130_fd_sc_hd__decap_3 PHY_5473 ();
 sky130_fd_sc_hd__decap_3 PHY_5474 ();
 sky130_fd_sc_hd__decap_3 PHY_5475 ();
 sky130_fd_sc_hd__decap_3 PHY_5476 ();
 sky130_fd_sc_hd__decap_3 PHY_5477 ();
 sky130_fd_sc_hd__decap_3 PHY_5478 ();
 sky130_fd_sc_hd__decap_3 PHY_5479 ();
 sky130_fd_sc_hd__decap_3 PHY_5480 ();
 sky130_fd_sc_hd__decap_3 PHY_5481 ();
 sky130_fd_sc_hd__decap_3 PHY_5482 ();
 sky130_fd_sc_hd__decap_3 PHY_5483 ();
 sky130_fd_sc_hd__decap_3 PHY_5484 ();
 sky130_fd_sc_hd__decap_3 PHY_5485 ();
 sky130_fd_sc_hd__decap_3 PHY_5486 ();
 sky130_fd_sc_hd__decap_3 PHY_5487 ();
 sky130_fd_sc_hd__decap_3 PHY_5488 ();
 sky130_fd_sc_hd__decap_3 PHY_5489 ();
 sky130_fd_sc_hd__decap_3 PHY_5490 ();
 sky130_fd_sc_hd__decap_3 PHY_5491 ();
 sky130_fd_sc_hd__decap_3 PHY_5492 ();
 sky130_fd_sc_hd__decap_3 PHY_5493 ();
 sky130_fd_sc_hd__decap_3 PHY_5494 ();
 sky130_fd_sc_hd__decap_3 PHY_5495 ();
 sky130_fd_sc_hd__decap_3 PHY_5496 ();
 sky130_fd_sc_hd__decap_3 PHY_5497 ();
 sky130_fd_sc_hd__decap_3 PHY_5498 ();
 sky130_fd_sc_hd__decap_3 PHY_5499 ();
 sky130_fd_sc_hd__decap_3 PHY_5500 ();
 sky130_fd_sc_hd__decap_3 PHY_5501 ();
 sky130_fd_sc_hd__decap_3 PHY_5502 ();
 sky130_fd_sc_hd__decap_3 PHY_5503 ();
 sky130_fd_sc_hd__decap_3 PHY_5504 ();
 sky130_fd_sc_hd__decap_3 PHY_5505 ();
 sky130_fd_sc_hd__decap_3 PHY_5506 ();
 sky130_fd_sc_hd__decap_3 PHY_5507 ();
 sky130_fd_sc_hd__decap_3 PHY_5508 ();
 sky130_fd_sc_hd__decap_3 PHY_5509 ();
 sky130_fd_sc_hd__decap_3 PHY_5510 ();
 sky130_fd_sc_hd__decap_3 PHY_5511 ();
 sky130_fd_sc_hd__decap_3 PHY_5512 ();
 sky130_fd_sc_hd__decap_3 PHY_5513 ();
 sky130_fd_sc_hd__decap_3 PHY_5514 ();
 sky130_fd_sc_hd__decap_3 PHY_5515 ();
 sky130_fd_sc_hd__decap_3 PHY_5516 ();
 sky130_fd_sc_hd__decap_3 PHY_5517 ();
 sky130_fd_sc_hd__decap_3 PHY_5518 ();
 sky130_fd_sc_hd__decap_3 PHY_5519 ();
 sky130_fd_sc_hd__decap_3 PHY_5520 ();
 sky130_fd_sc_hd__decap_3 PHY_5521 ();
 sky130_fd_sc_hd__decap_3 PHY_5522 ();
 sky130_fd_sc_hd__decap_3 PHY_5523 ();
 sky130_fd_sc_hd__decap_3 PHY_5524 ();
 sky130_fd_sc_hd__decap_3 PHY_5525 ();
 sky130_fd_sc_hd__decap_3 PHY_5526 ();
 sky130_fd_sc_hd__decap_3 PHY_5527 ();
 sky130_fd_sc_hd__decap_3 PHY_5528 ();
 sky130_fd_sc_hd__decap_3 PHY_5529 ();
 sky130_fd_sc_hd__decap_3 PHY_5530 ();
 sky130_fd_sc_hd__decap_3 PHY_5531 ();
 sky130_fd_sc_hd__decap_3 PHY_5532 ();
 sky130_fd_sc_hd__decap_3 PHY_5533 ();
 sky130_fd_sc_hd__decap_3 PHY_5534 ();
 sky130_fd_sc_hd__decap_3 PHY_5535 ();
 sky130_fd_sc_hd__decap_3 PHY_5536 ();
 sky130_fd_sc_hd__decap_3 PHY_5537 ();
 sky130_fd_sc_hd__decap_3 PHY_5538 ();
 sky130_fd_sc_hd__decap_3 PHY_5539 ();
 sky130_fd_sc_hd__decap_3 PHY_5540 ();
 sky130_fd_sc_hd__decap_3 PHY_5541 ();
 sky130_fd_sc_hd__decap_3 PHY_5542 ();
 sky130_fd_sc_hd__decap_3 PHY_5543 ();
 sky130_fd_sc_hd__decap_3 PHY_5544 ();
 sky130_fd_sc_hd__decap_3 PHY_5545 ();
 sky130_fd_sc_hd__decap_3 PHY_5546 ();
 sky130_fd_sc_hd__decap_3 PHY_5547 ();
 sky130_fd_sc_hd__decap_3 PHY_5548 ();
 sky130_fd_sc_hd__decap_3 PHY_5549 ();
 sky130_fd_sc_hd__decap_3 PHY_5550 ();
 sky130_fd_sc_hd__decap_3 PHY_5551 ();
 sky130_fd_sc_hd__decap_3 PHY_5552 ();
 sky130_fd_sc_hd__decap_3 PHY_5553 ();
 sky130_fd_sc_hd__decap_3 PHY_5554 ();
 sky130_fd_sc_hd__decap_3 PHY_5555 ();
 sky130_fd_sc_hd__decap_3 PHY_5556 ();
 sky130_fd_sc_hd__decap_3 PHY_5557 ();
 sky130_fd_sc_hd__decap_3 PHY_5558 ();
 sky130_fd_sc_hd__decap_3 PHY_5559 ();
 sky130_fd_sc_hd__decap_3 PHY_5560 ();
 sky130_fd_sc_hd__decap_3 PHY_5561 ();
 sky130_fd_sc_hd__decap_3 PHY_5562 ();
 sky130_fd_sc_hd__decap_3 PHY_5563 ();
 sky130_fd_sc_hd__decap_3 PHY_5564 ();
 sky130_fd_sc_hd__decap_3 PHY_5565 ();
 sky130_fd_sc_hd__decap_3 PHY_5566 ();
 sky130_fd_sc_hd__decap_3 PHY_5567 ();
 sky130_fd_sc_hd__decap_3 PHY_5568 ();
 sky130_fd_sc_hd__decap_3 PHY_5569 ();
 sky130_fd_sc_hd__decap_3 PHY_5570 ();
 sky130_fd_sc_hd__decap_3 PHY_5571 ();
 sky130_fd_sc_hd__decap_3 PHY_5572 ();
 sky130_fd_sc_hd__decap_3 PHY_5573 ();
 sky130_fd_sc_hd__decap_3 PHY_5574 ();
 sky130_fd_sc_hd__decap_3 PHY_5575 ();
 sky130_fd_sc_hd__decap_3 PHY_5576 ();
 sky130_fd_sc_hd__decap_3 PHY_5577 ();
 sky130_fd_sc_hd__decap_3 PHY_5578 ();
 sky130_fd_sc_hd__decap_3 PHY_5579 ();
 sky130_fd_sc_hd__decap_3 PHY_5580 ();
 sky130_fd_sc_hd__decap_3 PHY_5581 ();
 sky130_fd_sc_hd__decap_3 PHY_5582 ();
 sky130_fd_sc_hd__decap_3 PHY_5583 ();
 sky130_fd_sc_hd__decap_3 PHY_5584 ();
 sky130_fd_sc_hd__decap_3 PHY_5585 ();
 sky130_fd_sc_hd__decap_3 PHY_5586 ();
 sky130_fd_sc_hd__decap_3 PHY_5587 ();
 sky130_fd_sc_hd__decap_3 PHY_5588 ();
 sky130_fd_sc_hd__decap_3 PHY_5589 ();
 sky130_fd_sc_hd__decap_3 PHY_5590 ();
 sky130_fd_sc_hd__decap_3 PHY_5591 ();
 sky130_fd_sc_hd__decap_3 PHY_5592 ();
 sky130_fd_sc_hd__decap_3 PHY_5593 ();
 sky130_fd_sc_hd__decap_3 PHY_5594 ();
 sky130_fd_sc_hd__decap_3 PHY_5595 ();
 sky130_fd_sc_hd__decap_3 PHY_5596 ();
 sky130_fd_sc_hd__decap_3 PHY_5597 ();
 sky130_fd_sc_hd__decap_3 PHY_5598 ();
 sky130_fd_sc_hd__decap_3 PHY_5599 ();
 sky130_fd_sc_hd__decap_3 PHY_5600 ();
 sky130_fd_sc_hd__decap_3 PHY_5601 ();
 sky130_fd_sc_hd__decap_3 PHY_5602 ();
 sky130_fd_sc_hd__decap_3 PHY_5603 ();
 sky130_fd_sc_hd__decap_3 PHY_5604 ();
 sky130_fd_sc_hd__decap_3 PHY_5605 ();
 sky130_fd_sc_hd__decap_3 PHY_5606 ();
 sky130_fd_sc_hd__decap_3 PHY_5607 ();
 sky130_fd_sc_hd__decap_3 PHY_5608 ();
 sky130_fd_sc_hd__decap_3 PHY_5609 ();
 sky130_fd_sc_hd__decap_3 PHY_5610 ();
 sky130_fd_sc_hd__decap_3 PHY_5611 ();
 sky130_fd_sc_hd__decap_3 PHY_5612 ();
 sky130_fd_sc_hd__decap_3 PHY_5613 ();
 sky130_fd_sc_hd__decap_3 PHY_5614 ();
 sky130_fd_sc_hd__decap_3 PHY_5615 ();
 sky130_fd_sc_hd__decap_3 PHY_5616 ();
 sky130_fd_sc_hd__decap_3 PHY_5617 ();
 sky130_fd_sc_hd__decap_3 PHY_5618 ();
 sky130_fd_sc_hd__decap_3 PHY_5619 ();
 sky130_fd_sc_hd__decap_3 PHY_5620 ();
 sky130_fd_sc_hd__decap_3 PHY_5621 ();
 sky130_fd_sc_hd__decap_3 PHY_5622 ();
 sky130_fd_sc_hd__decap_3 PHY_5623 ();
 sky130_fd_sc_hd__decap_3 PHY_5624 ();
 sky130_fd_sc_hd__decap_3 PHY_5625 ();
 sky130_fd_sc_hd__decap_3 PHY_5626 ();
 sky130_fd_sc_hd__decap_3 PHY_5627 ();
 sky130_fd_sc_hd__decap_3 PHY_5628 ();
 sky130_fd_sc_hd__decap_3 PHY_5629 ();
 sky130_fd_sc_hd__decap_3 PHY_5630 ();
 sky130_fd_sc_hd__decap_3 PHY_5631 ();
 sky130_fd_sc_hd__decap_3 PHY_5632 ();
 sky130_fd_sc_hd__decap_3 PHY_5633 ();
 sky130_fd_sc_hd__decap_3 PHY_5634 ();
 sky130_fd_sc_hd__decap_3 PHY_5635 ();
 sky130_fd_sc_hd__decap_3 PHY_5636 ();
 sky130_fd_sc_hd__decap_3 PHY_5637 ();
 sky130_fd_sc_hd__decap_3 PHY_5638 ();
 sky130_fd_sc_hd__decap_3 PHY_5639 ();
 sky130_fd_sc_hd__decap_3 PHY_5640 ();
 sky130_fd_sc_hd__decap_3 PHY_5641 ();
 sky130_fd_sc_hd__decap_3 PHY_5642 ();
 sky130_fd_sc_hd__decap_3 PHY_5643 ();
 sky130_fd_sc_hd__decap_3 PHY_5644 ();
 sky130_fd_sc_hd__decap_3 PHY_5645 ();
 sky130_fd_sc_hd__decap_3 PHY_5646 ();
 sky130_fd_sc_hd__decap_3 PHY_5647 ();
 sky130_fd_sc_hd__decap_3 PHY_5648 ();
 sky130_fd_sc_hd__decap_3 PHY_5649 ();
 sky130_fd_sc_hd__decap_3 PHY_5650 ();
 sky130_fd_sc_hd__decap_3 PHY_5651 ();
 sky130_fd_sc_hd__decap_3 PHY_5652 ();
 sky130_fd_sc_hd__decap_3 PHY_5653 ();
 sky130_fd_sc_hd__decap_3 PHY_5654 ();
 sky130_fd_sc_hd__decap_3 PHY_5655 ();
 sky130_fd_sc_hd__decap_3 PHY_5656 ();
 sky130_fd_sc_hd__decap_3 PHY_5657 ();
 sky130_fd_sc_hd__decap_3 PHY_5658 ();
 sky130_fd_sc_hd__decap_3 PHY_5659 ();
 sky130_fd_sc_hd__decap_3 PHY_5660 ();
 sky130_fd_sc_hd__decap_3 PHY_5661 ();
 sky130_fd_sc_hd__decap_3 PHY_5662 ();
 sky130_fd_sc_hd__decap_3 PHY_5663 ();
 sky130_fd_sc_hd__decap_3 PHY_5664 ();
 sky130_fd_sc_hd__decap_3 PHY_5665 ();
 sky130_fd_sc_hd__decap_3 PHY_5666 ();
 sky130_fd_sc_hd__decap_3 PHY_5667 ();
 sky130_fd_sc_hd__decap_3 PHY_5668 ();
 sky130_fd_sc_hd__decap_3 PHY_5669 ();
 sky130_fd_sc_hd__decap_3 PHY_5670 ();
 sky130_fd_sc_hd__decap_3 PHY_5671 ();
 sky130_fd_sc_hd__decap_3 PHY_5672 ();
 sky130_fd_sc_hd__decap_3 PHY_5673 ();
 sky130_fd_sc_hd__decap_3 PHY_5674 ();
 sky130_fd_sc_hd__decap_3 PHY_5675 ();
 sky130_fd_sc_hd__decap_3 PHY_5676 ();
 sky130_fd_sc_hd__decap_3 PHY_5677 ();
 sky130_fd_sc_hd__decap_3 PHY_5678 ();
 sky130_fd_sc_hd__decap_3 PHY_5679 ();
 sky130_fd_sc_hd__decap_3 PHY_5680 ();
 sky130_fd_sc_hd__decap_3 PHY_5681 ();
 sky130_fd_sc_hd__decap_3 PHY_5682 ();
 sky130_fd_sc_hd__decap_3 PHY_5683 ();
 sky130_fd_sc_hd__decap_3 PHY_5684 ();
 sky130_fd_sc_hd__decap_3 PHY_5685 ();
 sky130_fd_sc_hd__decap_3 PHY_5686 ();
 sky130_fd_sc_hd__decap_3 PHY_5687 ();
 sky130_fd_sc_hd__decap_3 PHY_5688 ();
 sky130_fd_sc_hd__decap_3 PHY_5689 ();
 sky130_fd_sc_hd__decap_3 PHY_5690 ();
 sky130_fd_sc_hd__decap_3 PHY_5691 ();
 sky130_fd_sc_hd__decap_3 PHY_5692 ();
 sky130_fd_sc_hd__decap_3 PHY_5693 ();
 sky130_fd_sc_hd__decap_3 PHY_5694 ();
 sky130_fd_sc_hd__decap_3 PHY_5695 ();
 sky130_fd_sc_hd__decap_3 PHY_5696 ();
 sky130_fd_sc_hd__decap_3 PHY_5697 ();
 sky130_fd_sc_hd__decap_3 PHY_5698 ();
 sky130_fd_sc_hd__decap_3 PHY_5699 ();
 sky130_fd_sc_hd__decap_3 PHY_5700 ();
 sky130_fd_sc_hd__decap_3 PHY_5701 ();
 sky130_fd_sc_hd__decap_3 PHY_5702 ();
 sky130_fd_sc_hd__decap_3 PHY_5703 ();
 sky130_fd_sc_hd__decap_3 PHY_5704 ();
 sky130_fd_sc_hd__decap_3 PHY_5705 ();
 sky130_fd_sc_hd__decap_3 PHY_5706 ();
 sky130_fd_sc_hd__decap_3 PHY_5707 ();
 sky130_fd_sc_hd__decap_3 PHY_5708 ();
 sky130_fd_sc_hd__decap_3 PHY_5709 ();
 sky130_fd_sc_hd__decap_3 PHY_5710 ();
 sky130_fd_sc_hd__decap_3 PHY_5711 ();
 sky130_fd_sc_hd__decap_3 PHY_5712 ();
 sky130_fd_sc_hd__decap_3 PHY_5713 ();
 sky130_fd_sc_hd__decap_3 PHY_5714 ();
 sky130_fd_sc_hd__decap_3 PHY_5715 ();
 sky130_fd_sc_hd__decap_3 PHY_5716 ();
 sky130_fd_sc_hd__decap_3 PHY_5717 ();
 sky130_fd_sc_hd__decap_3 PHY_5718 ();
 sky130_fd_sc_hd__decap_3 PHY_5719 ();
 sky130_fd_sc_hd__decap_3 PHY_5720 ();
 sky130_fd_sc_hd__decap_3 PHY_5721 ();
 sky130_fd_sc_hd__decap_3 PHY_5722 ();
 sky130_fd_sc_hd__decap_3 PHY_5723 ();
 sky130_fd_sc_hd__decap_3 PHY_5724 ();
 sky130_fd_sc_hd__decap_3 PHY_5725 ();
 sky130_fd_sc_hd__decap_3 PHY_5726 ();
 sky130_fd_sc_hd__decap_3 PHY_5727 ();
 sky130_fd_sc_hd__decap_3 PHY_5728 ();
 sky130_fd_sc_hd__decap_3 PHY_5729 ();
 sky130_fd_sc_hd__decap_3 PHY_5730 ();
 sky130_fd_sc_hd__decap_3 PHY_5731 ();
 sky130_fd_sc_hd__decap_3 PHY_5732 ();
 sky130_fd_sc_hd__decap_3 PHY_5733 ();
 sky130_fd_sc_hd__decap_3 PHY_5734 ();
 sky130_fd_sc_hd__decap_3 PHY_5735 ();
 sky130_fd_sc_hd__decap_3 PHY_5736 ();
 sky130_fd_sc_hd__decap_3 PHY_5737 ();
 sky130_fd_sc_hd__decap_3 PHY_5738 ();
 sky130_fd_sc_hd__decap_3 PHY_5739 ();
 sky130_fd_sc_hd__decap_3 PHY_5740 ();
 sky130_fd_sc_hd__decap_3 PHY_5741 ();
 sky130_fd_sc_hd__decap_3 PHY_5742 ();
 sky130_fd_sc_hd__decap_3 PHY_5743 ();
 sky130_fd_sc_hd__decap_3 PHY_5744 ();
 sky130_fd_sc_hd__decap_3 PHY_5745 ();
 sky130_fd_sc_hd__decap_3 PHY_5746 ();
 sky130_fd_sc_hd__decap_3 PHY_5747 ();
 sky130_fd_sc_hd__decap_3 PHY_5748 ();
 sky130_fd_sc_hd__decap_3 PHY_5749 ();
 sky130_fd_sc_hd__decap_3 PHY_5750 ();
 sky130_fd_sc_hd__decap_3 PHY_5751 ();
 sky130_fd_sc_hd__decap_3 PHY_5752 ();
 sky130_fd_sc_hd__decap_3 PHY_5753 ();
 sky130_fd_sc_hd__decap_3 PHY_5754 ();
 sky130_fd_sc_hd__decap_3 PHY_5755 ();
 sky130_fd_sc_hd__decap_3 PHY_5756 ();
 sky130_fd_sc_hd__decap_3 PHY_5757 ();
 sky130_fd_sc_hd__decap_3 PHY_5758 ();
 sky130_fd_sc_hd__decap_3 PHY_5759 ();
 sky130_fd_sc_hd__decap_3 PHY_5760 ();
 sky130_fd_sc_hd__decap_3 PHY_5761 ();
 sky130_fd_sc_hd__decap_3 PHY_5762 ();
 sky130_fd_sc_hd__decap_3 PHY_5763 ();
 sky130_fd_sc_hd__decap_3 PHY_5764 ();
 sky130_fd_sc_hd__decap_3 PHY_5765 ();
 sky130_fd_sc_hd__decap_3 PHY_5766 ();
 sky130_fd_sc_hd__decap_3 PHY_5767 ();
 sky130_fd_sc_hd__decap_3 PHY_5768 ();
 sky130_fd_sc_hd__decap_3 PHY_5769 ();
 sky130_fd_sc_hd__decap_3 PHY_5770 ();
 sky130_fd_sc_hd__decap_3 PHY_5771 ();
 sky130_fd_sc_hd__decap_3 PHY_5772 ();
 sky130_fd_sc_hd__decap_3 PHY_5773 ();
 sky130_fd_sc_hd__decap_3 PHY_5774 ();
 sky130_fd_sc_hd__decap_3 PHY_5775 ();
 sky130_fd_sc_hd__decap_3 PHY_5776 ();
 sky130_fd_sc_hd__decap_3 PHY_5777 ();
 sky130_fd_sc_hd__decap_3 PHY_5778 ();
 sky130_fd_sc_hd__decap_3 PHY_5779 ();
 sky130_fd_sc_hd__decap_3 PHY_5780 ();
 sky130_fd_sc_hd__decap_3 PHY_5781 ();
 sky130_fd_sc_hd__decap_3 PHY_5782 ();
 sky130_fd_sc_hd__decap_3 PHY_5783 ();
 sky130_fd_sc_hd__decap_3 PHY_5784 ();
 sky130_fd_sc_hd__decap_3 PHY_5785 ();
 sky130_fd_sc_hd__decap_3 PHY_5786 ();
 sky130_fd_sc_hd__decap_3 PHY_5787 ();
 sky130_fd_sc_hd__decap_3 PHY_5788 ();
 sky130_fd_sc_hd__decap_3 PHY_5789 ();
 sky130_fd_sc_hd__decap_3 PHY_5790 ();
 sky130_fd_sc_hd__decap_3 PHY_5791 ();
 sky130_fd_sc_hd__decap_3 PHY_5792 ();
 sky130_fd_sc_hd__decap_3 PHY_5793 ();
 sky130_fd_sc_hd__decap_3 PHY_5794 ();
 sky130_fd_sc_hd__decap_3 PHY_5795 ();
 sky130_fd_sc_hd__decap_3 PHY_5796 ();
 sky130_fd_sc_hd__decap_3 PHY_5797 ();
 sky130_fd_sc_hd__decap_3 PHY_5798 ();
 sky130_fd_sc_hd__decap_3 PHY_5799 ();
 sky130_fd_sc_hd__decap_3 PHY_5800 ();
 sky130_fd_sc_hd__decap_3 PHY_5801 ();
 sky130_fd_sc_hd__decap_3 PHY_5802 ();
 sky130_fd_sc_hd__decap_3 PHY_5803 ();
 sky130_fd_sc_hd__decap_3 PHY_5804 ();
 sky130_fd_sc_hd__decap_3 PHY_5805 ();
 sky130_fd_sc_hd__decap_3 PHY_5806 ();
 sky130_fd_sc_hd__decap_3 PHY_5807 ();
 sky130_fd_sc_hd__decap_3 PHY_5808 ();
 sky130_fd_sc_hd__decap_3 PHY_5809 ();
 sky130_fd_sc_hd__decap_3 PHY_5810 ();
 sky130_fd_sc_hd__decap_3 PHY_5811 ();
 sky130_fd_sc_hd__decap_3 PHY_5812 ();
 sky130_fd_sc_hd__decap_3 PHY_5813 ();
 sky130_fd_sc_hd__decap_3 PHY_5814 ();
 sky130_fd_sc_hd__decap_3 PHY_5815 ();
 sky130_fd_sc_hd__decap_3 PHY_5816 ();
 sky130_fd_sc_hd__decap_3 PHY_5817 ();
 sky130_fd_sc_hd__decap_3 PHY_5818 ();
 sky130_fd_sc_hd__decap_3 PHY_5819 ();
 sky130_fd_sc_hd__decap_3 PHY_5820 ();
 sky130_fd_sc_hd__decap_3 PHY_5821 ();
 sky130_fd_sc_hd__decap_3 PHY_5822 ();
 sky130_fd_sc_hd__decap_3 PHY_5823 ();
 sky130_fd_sc_hd__decap_3 PHY_5824 ();
 sky130_fd_sc_hd__decap_3 PHY_5825 ();
 sky130_fd_sc_hd__decap_3 PHY_5826 ();
 sky130_fd_sc_hd__decap_3 PHY_5827 ();
 sky130_fd_sc_hd__decap_3 PHY_5828 ();
 sky130_fd_sc_hd__decap_3 PHY_5829 ();
 sky130_fd_sc_hd__decap_3 PHY_5830 ();
 sky130_fd_sc_hd__decap_3 PHY_5831 ();
 sky130_fd_sc_hd__decap_3 PHY_5832 ();
 sky130_fd_sc_hd__decap_3 PHY_5833 ();
 sky130_fd_sc_hd__decap_3 PHY_5834 ();
 sky130_fd_sc_hd__decap_3 PHY_5835 ();
 sky130_fd_sc_hd__decap_3 PHY_5836 ();
 sky130_fd_sc_hd__decap_3 PHY_5837 ();
 sky130_fd_sc_hd__decap_3 PHY_5838 ();
 sky130_fd_sc_hd__decap_3 PHY_5839 ();
 sky130_fd_sc_hd__decap_3 PHY_5840 ();
 sky130_fd_sc_hd__decap_3 PHY_5841 ();
 sky130_fd_sc_hd__decap_3 PHY_5842 ();
 sky130_fd_sc_hd__decap_3 PHY_5843 ();
 sky130_fd_sc_hd__decap_3 PHY_5844 ();
 sky130_fd_sc_hd__decap_3 PHY_5845 ();
 sky130_fd_sc_hd__decap_3 PHY_5846 ();
 sky130_fd_sc_hd__decap_3 PHY_5847 ();
 sky130_fd_sc_hd__decap_3 PHY_5848 ();
 sky130_fd_sc_hd__decap_3 PHY_5849 ();
 sky130_fd_sc_hd__decap_3 PHY_5850 ();
 sky130_fd_sc_hd__decap_3 PHY_5851 ();
 sky130_fd_sc_hd__decap_3 PHY_5852 ();
 sky130_fd_sc_hd__decap_3 PHY_5853 ();
 sky130_fd_sc_hd__decap_3 PHY_5854 ();
 sky130_fd_sc_hd__decap_3 PHY_5855 ();
 sky130_fd_sc_hd__decap_3 PHY_5856 ();
 sky130_fd_sc_hd__decap_3 PHY_5857 ();
 sky130_fd_sc_hd__decap_3 PHY_5858 ();
 sky130_fd_sc_hd__decap_3 PHY_5859 ();
 sky130_fd_sc_hd__decap_3 PHY_5860 ();
 sky130_fd_sc_hd__decap_3 PHY_5861 ();
 sky130_fd_sc_hd__decap_3 PHY_5862 ();
 sky130_fd_sc_hd__decap_3 PHY_5863 ();
 sky130_fd_sc_hd__decap_3 PHY_5864 ();
 sky130_fd_sc_hd__decap_3 PHY_5865 ();
 sky130_fd_sc_hd__decap_3 PHY_5866 ();
 sky130_fd_sc_hd__decap_3 PHY_5867 ();
 sky130_fd_sc_hd__decap_3 PHY_5868 ();
 sky130_fd_sc_hd__decap_3 PHY_5869 ();
 sky130_fd_sc_hd__decap_3 PHY_5870 ();
 sky130_fd_sc_hd__decap_3 PHY_5871 ();
 sky130_fd_sc_hd__decap_3 PHY_5872 ();
 sky130_fd_sc_hd__decap_3 PHY_5873 ();
 sky130_fd_sc_hd__decap_3 PHY_5874 ();
 sky130_fd_sc_hd__decap_3 PHY_5875 ();
 sky130_fd_sc_hd__decap_3 PHY_5876 ();
 sky130_fd_sc_hd__decap_3 PHY_5877 ();
 sky130_fd_sc_hd__decap_3 PHY_5878 ();
 sky130_fd_sc_hd__decap_3 PHY_5879 ();
 sky130_fd_sc_hd__decap_3 PHY_5880 ();
 sky130_fd_sc_hd__decap_3 PHY_5881 ();
 sky130_fd_sc_hd__decap_3 PHY_5882 ();
 sky130_fd_sc_hd__decap_3 PHY_5883 ();
 sky130_fd_sc_hd__decap_3 PHY_5884 ();
 sky130_fd_sc_hd__decap_3 PHY_5885 ();
 sky130_fd_sc_hd__decap_3 PHY_5886 ();
 sky130_fd_sc_hd__decap_3 PHY_5887 ();
 sky130_fd_sc_hd__decap_3 PHY_5888 ();
 sky130_fd_sc_hd__decap_3 PHY_5889 ();
 sky130_fd_sc_hd__decap_3 PHY_5890 ();
 sky130_fd_sc_hd__decap_3 PHY_5891 ();
 sky130_fd_sc_hd__decap_3 PHY_5892 ();
 sky130_fd_sc_hd__decap_3 PHY_5893 ();
 sky130_fd_sc_hd__decap_3 PHY_5894 ();
 sky130_fd_sc_hd__decap_3 PHY_5895 ();
 sky130_fd_sc_hd__decap_3 PHY_5896 ();
 sky130_fd_sc_hd__decap_3 PHY_5897 ();
 sky130_fd_sc_hd__decap_3 PHY_5898 ();
 sky130_fd_sc_hd__decap_3 PHY_5899 ();
 sky130_fd_sc_hd__decap_3 PHY_5900 ();
 sky130_fd_sc_hd__decap_3 PHY_5901 ();
 sky130_fd_sc_hd__decap_3 PHY_5902 ();
 sky130_fd_sc_hd__decap_3 PHY_5903 ();
 sky130_fd_sc_hd__decap_3 PHY_5904 ();
 sky130_fd_sc_hd__decap_3 PHY_5905 ();
 sky130_fd_sc_hd__decap_3 PHY_5906 ();
 sky130_fd_sc_hd__decap_3 PHY_5907 ();
 sky130_fd_sc_hd__decap_3 PHY_5908 ();
 sky130_fd_sc_hd__decap_3 PHY_5909 ();
 sky130_fd_sc_hd__decap_3 PHY_5910 ();
 sky130_fd_sc_hd__decap_3 PHY_5911 ();
 sky130_fd_sc_hd__decap_3 PHY_5912 ();
 sky130_fd_sc_hd__decap_3 PHY_5913 ();
 sky130_fd_sc_hd__decap_3 PHY_5914 ();
 sky130_fd_sc_hd__decap_3 PHY_5915 ();
 sky130_fd_sc_hd__decap_3 PHY_5916 ();
 sky130_fd_sc_hd__decap_3 PHY_5917 ();
 sky130_fd_sc_hd__decap_3 PHY_5918 ();
 sky130_fd_sc_hd__decap_3 PHY_5919 ();
 sky130_fd_sc_hd__decap_3 PHY_5920 ();
 sky130_fd_sc_hd__decap_3 PHY_5921 ();
 sky130_fd_sc_hd__decap_3 PHY_5922 ();
 sky130_fd_sc_hd__decap_3 PHY_5923 ();
 sky130_fd_sc_hd__decap_3 PHY_5924 ();
 sky130_fd_sc_hd__decap_3 PHY_5925 ();
 sky130_fd_sc_hd__decap_3 PHY_5926 ();
 sky130_fd_sc_hd__decap_3 PHY_5927 ();
 sky130_fd_sc_hd__decap_3 PHY_5928 ();
 sky130_fd_sc_hd__decap_3 PHY_5929 ();
 sky130_fd_sc_hd__decap_3 PHY_5930 ();
 sky130_fd_sc_hd__decap_3 PHY_5931 ();
 sky130_fd_sc_hd__decap_3 PHY_5932 ();
 sky130_fd_sc_hd__decap_3 PHY_5933 ();
 sky130_fd_sc_hd__decap_3 PHY_5934 ();
 sky130_fd_sc_hd__decap_3 PHY_5935 ();
 sky130_fd_sc_hd__decap_3 PHY_5936 ();
 sky130_fd_sc_hd__decap_3 PHY_5937 ();
 sky130_fd_sc_hd__decap_3 PHY_5938 ();
 sky130_fd_sc_hd__decap_3 PHY_5939 ();
 sky130_fd_sc_hd__decap_3 PHY_5940 ();
 sky130_fd_sc_hd__decap_3 PHY_5941 ();
 sky130_fd_sc_hd__decap_3 PHY_5942 ();
 sky130_fd_sc_hd__decap_3 PHY_5943 ();
 sky130_fd_sc_hd__decap_3 PHY_5944 ();
 sky130_fd_sc_hd__decap_3 PHY_5945 ();
 sky130_fd_sc_hd__decap_3 PHY_5946 ();
 sky130_fd_sc_hd__decap_3 PHY_5947 ();
 sky130_fd_sc_hd__decap_3 PHY_5948 ();
 sky130_fd_sc_hd__decap_3 PHY_5949 ();
 sky130_fd_sc_hd__decap_3 PHY_5950 ();
 sky130_fd_sc_hd__decap_3 PHY_5951 ();
 sky130_fd_sc_hd__decap_3 PHY_5952 ();
 sky130_fd_sc_hd__decap_3 PHY_5953 ();
 sky130_fd_sc_hd__decap_3 PHY_5954 ();
 sky130_fd_sc_hd__decap_3 PHY_5955 ();
 sky130_fd_sc_hd__decap_3 PHY_5956 ();
 sky130_fd_sc_hd__decap_3 PHY_5957 ();
 sky130_fd_sc_hd__decap_3 PHY_5958 ();
 sky130_fd_sc_hd__decap_3 PHY_5959 ();
 sky130_fd_sc_hd__decap_3 PHY_5960 ();
 sky130_fd_sc_hd__decap_3 PHY_5961 ();
 sky130_fd_sc_hd__decap_3 PHY_5962 ();
 sky130_fd_sc_hd__decap_3 PHY_5963 ();
 sky130_fd_sc_hd__decap_3 PHY_5964 ();
 sky130_fd_sc_hd__decap_3 PHY_5965 ();
 sky130_fd_sc_hd__decap_3 PHY_5966 ();
 sky130_fd_sc_hd__decap_3 PHY_5967 ();
 sky130_fd_sc_hd__decap_3 PHY_5968 ();
 sky130_fd_sc_hd__decap_3 PHY_5969 ();
 sky130_fd_sc_hd__decap_3 PHY_5970 ();
 sky130_fd_sc_hd__decap_3 PHY_5971 ();
 sky130_fd_sc_hd__decap_3 PHY_5972 ();
 sky130_fd_sc_hd__decap_3 PHY_5973 ();
 sky130_fd_sc_hd__decap_3 PHY_5974 ();
 sky130_fd_sc_hd__decap_3 PHY_5975 ();
 sky130_fd_sc_hd__decap_3 PHY_5976 ();
 sky130_fd_sc_hd__decap_3 PHY_5977 ();
 sky130_fd_sc_hd__decap_3 PHY_5978 ();
 sky130_fd_sc_hd__decap_3 PHY_5979 ();
 sky130_fd_sc_hd__decap_3 PHY_5980 ();
 sky130_fd_sc_hd__decap_3 PHY_5981 ();
 sky130_fd_sc_hd__decap_3 PHY_5982 ();
 sky130_fd_sc_hd__decap_3 PHY_5983 ();
 sky130_fd_sc_hd__decap_3 PHY_5984 ();
 sky130_fd_sc_hd__decap_3 PHY_5985 ();
 sky130_fd_sc_hd__decap_3 PHY_5986 ();
 sky130_fd_sc_hd__decap_3 PHY_5987 ();
 sky130_fd_sc_hd__decap_3 PHY_5988 ();
 sky130_fd_sc_hd__decap_3 PHY_5989 ();
 sky130_fd_sc_hd__decap_3 PHY_5990 ();
 sky130_fd_sc_hd__decap_3 PHY_5991 ();
 sky130_fd_sc_hd__decap_3 PHY_5992 ();
 sky130_fd_sc_hd__decap_3 PHY_5993 ();
 sky130_fd_sc_hd__decap_3 PHY_5994 ();
 sky130_fd_sc_hd__decap_3 PHY_5995 ();
 sky130_fd_sc_hd__decap_3 PHY_5996 ();
 sky130_fd_sc_hd__decap_3 PHY_5997 ();
 sky130_fd_sc_hd__decap_3 PHY_5998 ();
 sky130_fd_sc_hd__decap_3 PHY_5999 ();
 sky130_fd_sc_hd__decap_3 PHY_6000 ();
 sky130_fd_sc_hd__decap_3 PHY_6001 ();
 sky130_fd_sc_hd__decap_3 PHY_6002 ();
 sky130_fd_sc_hd__decap_3 PHY_6003 ();
 sky130_fd_sc_hd__decap_3 PHY_6004 ();
 sky130_fd_sc_hd__decap_3 PHY_6005 ();
 sky130_fd_sc_hd__decap_3 PHY_6006 ();
 sky130_fd_sc_hd__decap_3 PHY_6007 ();
 sky130_fd_sc_hd__decap_3 PHY_6008 ();
 sky130_fd_sc_hd__decap_3 PHY_6009 ();
 sky130_fd_sc_hd__decap_3 PHY_6010 ();
 sky130_fd_sc_hd__decap_3 PHY_6011 ();
 sky130_fd_sc_hd__decap_3 PHY_6012 ();
 sky130_fd_sc_hd__decap_3 PHY_6013 ();
 sky130_fd_sc_hd__decap_3 PHY_6014 ();
 sky130_fd_sc_hd__decap_3 PHY_6015 ();
 sky130_fd_sc_hd__decap_3 PHY_6016 ();
 sky130_fd_sc_hd__decap_3 PHY_6017 ();
 sky130_fd_sc_hd__decap_3 PHY_6018 ();
 sky130_fd_sc_hd__decap_3 PHY_6019 ();
 sky130_fd_sc_hd__decap_3 PHY_6020 ();
 sky130_fd_sc_hd__decap_3 PHY_6021 ();
 sky130_fd_sc_hd__decap_3 PHY_6022 ();
 sky130_fd_sc_hd__decap_3 PHY_6023 ();
 sky130_fd_sc_hd__decap_3 PHY_6024 ();
 sky130_fd_sc_hd__decap_3 PHY_6025 ();
 sky130_fd_sc_hd__decap_3 PHY_6026 ();
 sky130_fd_sc_hd__decap_3 PHY_6027 ();
 sky130_fd_sc_hd__decap_3 PHY_6028 ();
 sky130_fd_sc_hd__decap_3 PHY_6029 ();
 sky130_fd_sc_hd__decap_3 PHY_6030 ();
 sky130_fd_sc_hd__decap_3 PHY_6031 ();
 sky130_fd_sc_hd__decap_3 PHY_6032 ();
 sky130_fd_sc_hd__decap_3 PHY_6033 ();
 sky130_fd_sc_hd__decap_3 PHY_6034 ();
 sky130_fd_sc_hd__decap_3 PHY_6035 ();
 sky130_fd_sc_hd__decap_3 PHY_6036 ();
 sky130_fd_sc_hd__decap_3 PHY_6037 ();
 sky130_fd_sc_hd__decap_3 PHY_6038 ();
 sky130_fd_sc_hd__decap_3 PHY_6039 ();
 sky130_fd_sc_hd__decap_3 PHY_6040 ();
 sky130_fd_sc_hd__decap_3 PHY_6041 ();
 sky130_fd_sc_hd__decap_3 PHY_6042 ();
 sky130_fd_sc_hd__decap_3 PHY_6043 ();
 sky130_fd_sc_hd__decap_3 PHY_6044 ();
 sky130_fd_sc_hd__decap_3 PHY_6045 ();
 sky130_fd_sc_hd__decap_3 PHY_6046 ();
 sky130_fd_sc_hd__decap_3 PHY_6047 ();
 sky130_fd_sc_hd__decap_3 PHY_6048 ();
 sky130_fd_sc_hd__decap_3 PHY_6049 ();
 sky130_fd_sc_hd__decap_3 PHY_6050 ();
 sky130_fd_sc_hd__decap_3 PHY_6051 ();
 sky130_fd_sc_hd__decap_3 PHY_6052 ();
 sky130_fd_sc_hd__decap_3 PHY_6053 ();
 sky130_fd_sc_hd__decap_3 PHY_6054 ();
 sky130_fd_sc_hd__decap_3 PHY_6055 ();
 sky130_fd_sc_hd__decap_3 PHY_6056 ();
 sky130_fd_sc_hd__decap_3 PHY_6057 ();
 sky130_fd_sc_hd__decap_3 PHY_6058 ();
 sky130_fd_sc_hd__decap_3 PHY_6059 ();
 sky130_fd_sc_hd__decap_3 PHY_6060 ();
 sky130_fd_sc_hd__decap_3 PHY_6061 ();
 sky130_fd_sc_hd__decap_3 PHY_6062 ();
 sky130_fd_sc_hd__decap_3 PHY_6063 ();
 sky130_fd_sc_hd__decap_3 PHY_6064 ();
 sky130_fd_sc_hd__decap_3 PHY_6065 ();
 sky130_fd_sc_hd__decap_3 PHY_6066 ();
 sky130_fd_sc_hd__decap_3 PHY_6067 ();
 sky130_fd_sc_hd__decap_3 PHY_6068 ();
 sky130_fd_sc_hd__decap_3 PHY_6069 ();
 sky130_fd_sc_hd__decap_3 PHY_6070 ();
 sky130_fd_sc_hd__decap_3 PHY_6071 ();
 sky130_fd_sc_hd__decap_3 PHY_6072 ();
 sky130_fd_sc_hd__decap_3 PHY_6073 ();
 sky130_fd_sc_hd__decap_3 PHY_6074 ();
 sky130_fd_sc_hd__decap_3 PHY_6075 ();
 sky130_fd_sc_hd__decap_3 PHY_6076 ();
 sky130_fd_sc_hd__decap_3 PHY_6077 ();
 sky130_fd_sc_hd__decap_3 PHY_6078 ();
 sky130_fd_sc_hd__decap_3 PHY_6079 ();
 sky130_fd_sc_hd__decap_3 PHY_6080 ();
 sky130_fd_sc_hd__decap_3 PHY_6081 ();
 sky130_fd_sc_hd__decap_3 PHY_6082 ();
 sky130_fd_sc_hd__decap_3 PHY_6083 ();
 sky130_fd_sc_hd__decap_3 PHY_6084 ();
 sky130_fd_sc_hd__decap_3 PHY_6085 ();
 sky130_fd_sc_hd__decap_3 PHY_6086 ();
 sky130_fd_sc_hd__decap_3 PHY_6087 ();
 sky130_fd_sc_hd__decap_3 PHY_6088 ();
 sky130_fd_sc_hd__decap_3 PHY_6089 ();
 sky130_fd_sc_hd__decap_3 PHY_6090 ();
 sky130_fd_sc_hd__decap_3 PHY_6091 ();
 sky130_fd_sc_hd__decap_3 PHY_6092 ();
 sky130_fd_sc_hd__decap_3 PHY_6093 ();
 sky130_fd_sc_hd__decap_3 PHY_6094 ();
 sky130_fd_sc_hd__decap_3 PHY_6095 ();
 sky130_fd_sc_hd__decap_3 PHY_6096 ();
 sky130_fd_sc_hd__decap_3 PHY_6097 ();
 sky130_fd_sc_hd__decap_3 PHY_6098 ();
 sky130_fd_sc_hd__decap_3 PHY_6099 ();
 sky130_fd_sc_hd__decap_3 PHY_6100 ();
 sky130_fd_sc_hd__decap_3 PHY_6101 ();
 sky130_fd_sc_hd__decap_3 PHY_6102 ();
 sky130_fd_sc_hd__decap_3 PHY_6103 ();
 sky130_fd_sc_hd__decap_3 PHY_6104 ();
 sky130_fd_sc_hd__decap_3 PHY_6105 ();
 sky130_fd_sc_hd__decap_3 PHY_6106 ();
 sky130_fd_sc_hd__decap_3 PHY_6107 ();
 sky130_fd_sc_hd__decap_3 PHY_6108 ();
 sky130_fd_sc_hd__decap_3 PHY_6109 ();
 sky130_fd_sc_hd__decap_3 PHY_6110 ();
 sky130_fd_sc_hd__decap_3 PHY_6111 ();
 sky130_fd_sc_hd__decap_3 PHY_6112 ();
 sky130_fd_sc_hd__decap_3 PHY_6113 ();
 sky130_fd_sc_hd__decap_3 PHY_6114 ();
 sky130_fd_sc_hd__decap_3 PHY_6115 ();
 sky130_fd_sc_hd__decap_3 PHY_6116 ();
 sky130_fd_sc_hd__decap_3 PHY_6117 ();
 sky130_fd_sc_hd__decap_3 PHY_6118 ();
 sky130_fd_sc_hd__decap_3 PHY_6119 ();
 sky130_fd_sc_hd__decap_3 PHY_6120 ();
 sky130_fd_sc_hd__decap_3 PHY_6121 ();
 sky130_fd_sc_hd__decap_3 PHY_6122 ();
 sky130_fd_sc_hd__decap_3 PHY_6123 ();
 sky130_fd_sc_hd__decap_3 PHY_6124 ();
 sky130_fd_sc_hd__decap_3 PHY_6125 ();
 sky130_fd_sc_hd__decap_3 PHY_6126 ();
 sky130_fd_sc_hd__decap_3 PHY_6127 ();
 sky130_fd_sc_hd__decap_3 PHY_6128 ();
 sky130_fd_sc_hd__decap_3 PHY_6129 ();
 sky130_fd_sc_hd__decap_3 PHY_6130 ();
 sky130_fd_sc_hd__decap_3 PHY_6131 ();
 sky130_fd_sc_hd__decap_3 PHY_6132 ();
 sky130_fd_sc_hd__decap_3 PHY_6133 ();
 sky130_fd_sc_hd__decap_3 PHY_6134 ();
 sky130_fd_sc_hd__decap_3 PHY_6135 ();
 sky130_fd_sc_hd__decap_3 PHY_6136 ();
 sky130_fd_sc_hd__decap_3 PHY_6137 ();
 sky130_fd_sc_hd__decap_3 PHY_6138 ();
 sky130_fd_sc_hd__decap_3 PHY_6139 ();
 sky130_fd_sc_hd__decap_3 PHY_6140 ();
 sky130_fd_sc_hd__decap_3 PHY_6141 ();
 sky130_fd_sc_hd__decap_3 PHY_6142 ();
 sky130_fd_sc_hd__decap_3 PHY_6143 ();
 sky130_fd_sc_hd__decap_3 PHY_6144 ();
 sky130_fd_sc_hd__decap_3 PHY_6145 ();
 sky130_fd_sc_hd__decap_3 PHY_6146 ();
 sky130_fd_sc_hd__decap_3 PHY_6147 ();
 sky130_fd_sc_hd__decap_3 PHY_6148 ();
 sky130_fd_sc_hd__decap_3 PHY_6149 ();
 sky130_fd_sc_hd__decap_3 PHY_6150 ();
 sky130_fd_sc_hd__decap_3 PHY_6151 ();
 sky130_fd_sc_hd__decap_3 PHY_6152 ();
 sky130_fd_sc_hd__decap_3 PHY_6153 ();
 sky130_fd_sc_hd__decap_3 PHY_6154 ();
 sky130_fd_sc_hd__decap_3 PHY_6155 ();
 sky130_fd_sc_hd__decap_3 PHY_6156 ();
 sky130_fd_sc_hd__decap_3 PHY_6157 ();
 sky130_fd_sc_hd__decap_3 PHY_6158 ();
 sky130_fd_sc_hd__decap_3 PHY_6159 ();
 sky130_fd_sc_hd__decap_3 PHY_6160 ();
 sky130_fd_sc_hd__decap_3 PHY_6161 ();
 sky130_fd_sc_hd__decap_3 PHY_6162 ();
 sky130_fd_sc_hd__decap_3 PHY_6163 ();
 sky130_fd_sc_hd__decap_3 PHY_6164 ();
 sky130_fd_sc_hd__decap_3 PHY_6165 ();
 sky130_fd_sc_hd__decap_3 PHY_6166 ();
 sky130_fd_sc_hd__decap_3 PHY_6167 ();
 sky130_fd_sc_hd__decap_3 PHY_6168 ();
 sky130_fd_sc_hd__decap_3 PHY_6169 ();
 sky130_fd_sc_hd__decap_3 PHY_6170 ();
 sky130_fd_sc_hd__decap_3 PHY_6171 ();
 sky130_fd_sc_hd__decap_3 PHY_6172 ();
 sky130_fd_sc_hd__decap_3 PHY_6173 ();
 sky130_fd_sc_hd__decap_3 PHY_6174 ();
 sky130_fd_sc_hd__decap_3 PHY_6175 ();
 sky130_fd_sc_hd__decap_3 PHY_6176 ();
 sky130_fd_sc_hd__decap_3 PHY_6177 ();
 sky130_fd_sc_hd__decap_3 PHY_6178 ();
 sky130_fd_sc_hd__decap_3 PHY_6179 ();
 sky130_fd_sc_hd__decap_3 PHY_6180 ();
 sky130_fd_sc_hd__decap_3 PHY_6181 ();
 sky130_fd_sc_hd__decap_3 PHY_6182 ();
 sky130_fd_sc_hd__decap_3 PHY_6183 ();
 sky130_fd_sc_hd__decap_3 PHY_6184 ();
 sky130_fd_sc_hd__decap_3 PHY_6185 ();
 sky130_fd_sc_hd__decap_3 PHY_6186 ();
 sky130_fd_sc_hd__decap_3 PHY_6187 ();
 sky130_fd_sc_hd__decap_3 PHY_6188 ();
 sky130_fd_sc_hd__decap_3 PHY_6189 ();
 sky130_fd_sc_hd__decap_3 PHY_6190 ();
 sky130_fd_sc_hd__decap_3 PHY_6191 ();
 sky130_fd_sc_hd__decap_3 PHY_6192 ();
 sky130_fd_sc_hd__decap_3 PHY_6193 ();
 sky130_fd_sc_hd__decap_3 PHY_6194 ();
 sky130_fd_sc_hd__decap_3 PHY_6195 ();
 sky130_fd_sc_hd__decap_3 PHY_6196 ();
 sky130_fd_sc_hd__decap_3 PHY_6197 ();
 sky130_fd_sc_hd__decap_3 PHY_6198 ();
 sky130_fd_sc_hd__decap_3 PHY_6199 ();
 sky130_fd_sc_hd__decap_3 PHY_6200 ();
 sky130_fd_sc_hd__decap_3 PHY_6201 ();
 sky130_fd_sc_hd__decap_3 PHY_6202 ();
 sky130_fd_sc_hd__decap_3 PHY_6203 ();
 sky130_fd_sc_hd__decap_3 PHY_6204 ();
 sky130_fd_sc_hd__decap_3 PHY_6205 ();
 sky130_fd_sc_hd__decap_3 PHY_6206 ();
 sky130_fd_sc_hd__decap_3 PHY_6207 ();
 sky130_fd_sc_hd__decap_3 PHY_6208 ();
 sky130_fd_sc_hd__decap_3 PHY_6209 ();
 sky130_fd_sc_hd__decap_3 PHY_6210 ();
 sky130_fd_sc_hd__decap_3 PHY_6211 ();
 sky130_fd_sc_hd__decap_3 PHY_6212 ();
 sky130_fd_sc_hd__decap_3 PHY_6213 ();
 sky130_fd_sc_hd__decap_3 PHY_6214 ();
 sky130_fd_sc_hd__decap_3 PHY_6215 ();
 sky130_fd_sc_hd__decap_3 PHY_6216 ();
 sky130_fd_sc_hd__decap_3 PHY_6217 ();
 sky130_fd_sc_hd__decap_3 PHY_6218 ();
 sky130_fd_sc_hd__decap_3 PHY_6219 ();
 sky130_fd_sc_hd__decap_3 PHY_6220 ();
 sky130_fd_sc_hd__decap_3 PHY_6221 ();
 sky130_fd_sc_hd__decap_3 PHY_6222 ();
 sky130_fd_sc_hd__decap_3 PHY_6223 ();
 sky130_fd_sc_hd__decap_3 PHY_6224 ();
 sky130_fd_sc_hd__decap_3 PHY_6225 ();
 sky130_fd_sc_hd__decap_3 PHY_6226 ();
 sky130_fd_sc_hd__decap_3 PHY_6227 ();
 sky130_fd_sc_hd__decap_3 PHY_6228 ();
 sky130_fd_sc_hd__decap_3 PHY_6229 ();
 sky130_fd_sc_hd__decap_3 PHY_6230 ();
 sky130_fd_sc_hd__decap_3 PHY_6231 ();
 sky130_fd_sc_hd__decap_3 PHY_6232 ();
 sky130_fd_sc_hd__decap_3 PHY_6233 ();
 sky130_fd_sc_hd__decap_3 PHY_6234 ();
 sky130_fd_sc_hd__decap_3 PHY_6235 ();
 sky130_fd_sc_hd__decap_3 PHY_6236 ();
 sky130_fd_sc_hd__decap_3 PHY_6237 ();
 sky130_fd_sc_hd__decap_3 PHY_6238 ();
 sky130_fd_sc_hd__decap_3 PHY_6239 ();
 sky130_fd_sc_hd__decap_3 PHY_6240 ();
 sky130_fd_sc_hd__decap_3 PHY_6241 ();
 sky130_fd_sc_hd__decap_3 PHY_6242 ();
 sky130_fd_sc_hd__decap_3 PHY_6243 ();
 sky130_fd_sc_hd__decap_3 PHY_6244 ();
 sky130_fd_sc_hd__decap_3 PHY_6245 ();
 sky130_fd_sc_hd__decap_3 PHY_6246 ();
 sky130_fd_sc_hd__decap_3 PHY_6247 ();
 sky130_fd_sc_hd__decap_3 PHY_6248 ();
 sky130_fd_sc_hd__decap_3 PHY_6249 ();
 sky130_fd_sc_hd__decap_3 PHY_6250 ();
 sky130_fd_sc_hd__decap_3 PHY_6251 ();
 sky130_fd_sc_hd__decap_3 PHY_6252 ();
 sky130_fd_sc_hd__decap_3 PHY_6253 ();
 sky130_fd_sc_hd__decap_3 PHY_6254 ();
 sky130_fd_sc_hd__decap_3 PHY_6255 ();
 sky130_fd_sc_hd__decap_3 PHY_6256 ();
 sky130_fd_sc_hd__decap_3 PHY_6257 ();
 sky130_fd_sc_hd__decap_3 PHY_6258 ();
 sky130_fd_sc_hd__decap_3 PHY_6259 ();
 sky130_fd_sc_hd__decap_3 PHY_6260 ();
 sky130_fd_sc_hd__decap_3 PHY_6261 ();
 sky130_fd_sc_hd__decap_3 PHY_6262 ();
 sky130_fd_sc_hd__decap_3 PHY_6263 ();
 sky130_fd_sc_hd__decap_3 PHY_6264 ();
 sky130_fd_sc_hd__decap_3 PHY_6265 ();
 sky130_fd_sc_hd__decap_3 PHY_6266 ();
 sky130_fd_sc_hd__decap_3 PHY_6267 ();
 sky130_fd_sc_hd__decap_3 PHY_6268 ();
 sky130_fd_sc_hd__decap_3 PHY_6269 ();
 sky130_fd_sc_hd__decap_3 PHY_6270 ();
 sky130_fd_sc_hd__decap_3 PHY_6271 ();
 sky130_fd_sc_hd__decap_3 PHY_6272 ();
 sky130_fd_sc_hd__decap_3 PHY_6273 ();
 sky130_fd_sc_hd__decap_3 PHY_6274 ();
 sky130_fd_sc_hd__decap_3 PHY_6275 ();
 sky130_fd_sc_hd__decap_3 PHY_6276 ();
 sky130_fd_sc_hd__decap_3 PHY_6277 ();
 sky130_fd_sc_hd__decap_3 PHY_6278 ();
 sky130_fd_sc_hd__decap_3 PHY_6279 ();
 sky130_fd_sc_hd__decap_3 PHY_6280 ();
 sky130_fd_sc_hd__decap_3 PHY_6281 ();
 sky130_fd_sc_hd__decap_3 PHY_6282 ();
 sky130_fd_sc_hd__decap_3 PHY_6283 ();
 sky130_fd_sc_hd__decap_3 PHY_6284 ();
 sky130_fd_sc_hd__decap_3 PHY_6285 ();
 sky130_fd_sc_hd__decap_3 PHY_6286 ();
 sky130_fd_sc_hd__decap_3 PHY_6287 ();
 sky130_fd_sc_hd__decap_3 PHY_6288 ();
 sky130_fd_sc_hd__decap_3 PHY_6289 ();
 sky130_fd_sc_hd__decap_3 PHY_6290 ();
 sky130_fd_sc_hd__decap_3 PHY_6291 ();
 sky130_fd_sc_hd__decap_3 PHY_6292 ();
 sky130_fd_sc_hd__decap_3 PHY_6293 ();
 sky130_fd_sc_hd__decap_3 PHY_6294 ();
 sky130_fd_sc_hd__decap_3 PHY_6295 ();
 sky130_fd_sc_hd__decap_3 PHY_6296 ();
 sky130_fd_sc_hd__decap_3 PHY_6297 ();
 sky130_fd_sc_hd__decap_3 PHY_6298 ();
 sky130_fd_sc_hd__decap_3 PHY_6299 ();
 sky130_fd_sc_hd__decap_3 PHY_6300 ();
 sky130_fd_sc_hd__decap_3 PHY_6301 ();
 sky130_fd_sc_hd__decap_3 PHY_6302 ();
 sky130_fd_sc_hd__decap_3 PHY_6303 ();
 sky130_fd_sc_hd__decap_3 PHY_6304 ();
 sky130_fd_sc_hd__decap_3 PHY_6305 ();
 sky130_fd_sc_hd__decap_3 PHY_6306 ();
 sky130_fd_sc_hd__decap_3 PHY_6307 ();
 sky130_fd_sc_hd__decap_3 PHY_6308 ();
 sky130_fd_sc_hd__decap_3 PHY_6309 ();
 sky130_fd_sc_hd__decap_3 PHY_6310 ();
 sky130_fd_sc_hd__decap_3 PHY_6311 ();
 sky130_fd_sc_hd__decap_3 PHY_6312 ();
 sky130_fd_sc_hd__decap_3 PHY_6313 ();
 sky130_fd_sc_hd__decap_3 PHY_6314 ();
 sky130_fd_sc_hd__decap_3 PHY_6315 ();
 sky130_fd_sc_hd__decap_3 PHY_6316 ();
 sky130_fd_sc_hd__decap_3 PHY_6317 ();
 sky130_fd_sc_hd__decap_3 PHY_6318 ();
 sky130_fd_sc_hd__decap_3 PHY_6319 ();
 sky130_fd_sc_hd__decap_3 PHY_6320 ();
 sky130_fd_sc_hd__decap_3 PHY_6321 ();
 sky130_fd_sc_hd__decap_3 PHY_6322 ();
 sky130_fd_sc_hd__decap_3 PHY_6323 ();
 sky130_fd_sc_hd__decap_3 PHY_6324 ();
 sky130_fd_sc_hd__decap_3 PHY_6325 ();
 sky130_fd_sc_hd__decap_3 PHY_6326 ();
 sky130_fd_sc_hd__decap_3 PHY_6327 ();
 sky130_fd_sc_hd__decap_3 PHY_6328 ();
 sky130_fd_sc_hd__decap_3 PHY_6329 ();
 sky130_fd_sc_hd__decap_3 PHY_6330 ();
 sky130_fd_sc_hd__decap_3 PHY_6331 ();
 sky130_fd_sc_hd__decap_3 PHY_6332 ();
 sky130_fd_sc_hd__decap_3 PHY_6333 ();
 sky130_fd_sc_hd__decap_3 PHY_6334 ();
 sky130_fd_sc_hd__decap_3 PHY_6335 ();
 sky130_fd_sc_hd__decap_3 PHY_6336 ();
 sky130_fd_sc_hd__decap_3 PHY_6337 ();
 sky130_fd_sc_hd__decap_3 PHY_6338 ();
 sky130_fd_sc_hd__decap_3 PHY_6339 ();
 sky130_fd_sc_hd__decap_3 PHY_6340 ();
 sky130_fd_sc_hd__decap_3 PHY_6341 ();
 sky130_fd_sc_hd__decap_3 PHY_6342 ();
 sky130_fd_sc_hd__decap_3 PHY_6343 ();
 sky130_fd_sc_hd__decap_3 PHY_6344 ();
 sky130_fd_sc_hd__decap_3 PHY_6345 ();
 sky130_fd_sc_hd__decap_3 PHY_6346 ();
 sky130_fd_sc_hd__decap_3 PHY_6347 ();
 sky130_fd_sc_hd__decap_3 PHY_6348 ();
 sky130_fd_sc_hd__decap_3 PHY_6349 ();
 sky130_fd_sc_hd__decap_3 PHY_6350 ();
 sky130_fd_sc_hd__decap_3 PHY_6351 ();
 sky130_fd_sc_hd__decap_3 PHY_6352 ();
 sky130_fd_sc_hd__decap_3 PHY_6353 ();
 sky130_fd_sc_hd__decap_3 PHY_6354 ();
 sky130_fd_sc_hd__decap_3 PHY_6355 ();
 sky130_fd_sc_hd__decap_3 PHY_6356 ();
 sky130_fd_sc_hd__decap_3 PHY_6357 ();
 sky130_fd_sc_hd__decap_3 PHY_6358 ();
 sky130_fd_sc_hd__decap_3 PHY_6359 ();
 sky130_fd_sc_hd__decap_3 PHY_6360 ();
 sky130_fd_sc_hd__decap_3 PHY_6361 ();
 sky130_fd_sc_hd__decap_3 PHY_6362 ();
 sky130_fd_sc_hd__decap_3 PHY_6363 ();
 sky130_fd_sc_hd__decap_3 PHY_6364 ();
 sky130_fd_sc_hd__decap_3 PHY_6365 ();
 sky130_fd_sc_hd__decap_3 PHY_6366 ();
 sky130_fd_sc_hd__decap_3 PHY_6367 ();
 sky130_fd_sc_hd__decap_3 PHY_6368 ();
 sky130_fd_sc_hd__decap_3 PHY_6369 ();
 sky130_fd_sc_hd__decap_3 PHY_6370 ();
 sky130_fd_sc_hd__decap_3 PHY_6371 ();
 sky130_fd_sc_hd__decap_3 PHY_6372 ();
 sky130_fd_sc_hd__decap_3 PHY_6373 ();
 sky130_fd_sc_hd__decap_3 PHY_6374 ();
 sky130_fd_sc_hd__decap_3 PHY_6375 ();
 sky130_fd_sc_hd__decap_3 PHY_6376 ();
 sky130_fd_sc_hd__decap_3 PHY_6377 ();
 sky130_fd_sc_hd__decap_3 PHY_6378 ();
 sky130_fd_sc_hd__decap_3 PHY_6379 ();
 sky130_fd_sc_hd__decap_3 PHY_6380 ();
 sky130_fd_sc_hd__decap_3 PHY_6381 ();
 sky130_fd_sc_hd__decap_3 PHY_6382 ();
 sky130_fd_sc_hd__decap_3 PHY_6383 ();
 sky130_fd_sc_hd__decap_3 PHY_6384 ();
 sky130_fd_sc_hd__decap_3 PHY_6385 ();
 sky130_fd_sc_hd__decap_3 PHY_6386 ();
 sky130_fd_sc_hd__decap_3 PHY_6387 ();
 sky130_fd_sc_hd__decap_3 PHY_6388 ();
 sky130_fd_sc_hd__decap_3 PHY_6389 ();
 sky130_fd_sc_hd__decap_3 PHY_6390 ();
 sky130_fd_sc_hd__decap_3 PHY_6391 ();
 sky130_fd_sc_hd__decap_3 PHY_6392 ();
 sky130_fd_sc_hd__decap_3 PHY_6393 ();
 sky130_fd_sc_hd__decap_3 PHY_6394 ();
 sky130_fd_sc_hd__decap_3 PHY_6395 ();
 sky130_fd_sc_hd__decap_3 PHY_6396 ();
 sky130_fd_sc_hd__decap_3 PHY_6397 ();
 sky130_fd_sc_hd__decap_3 PHY_6398 ();
 sky130_fd_sc_hd__decap_3 PHY_6399 ();
 sky130_fd_sc_hd__decap_3 PHY_6400 ();
 sky130_fd_sc_hd__decap_3 PHY_6401 ();
 sky130_fd_sc_hd__decap_3 PHY_6402 ();
 sky130_fd_sc_hd__decap_3 PHY_6403 ();
 sky130_fd_sc_hd__decap_3 PHY_6404 ();
 sky130_fd_sc_hd__decap_3 PHY_6405 ();
 sky130_fd_sc_hd__decap_3 PHY_6406 ();
 sky130_fd_sc_hd__decap_3 PHY_6407 ();
 sky130_fd_sc_hd__decap_3 PHY_6408 ();
 sky130_fd_sc_hd__decap_3 PHY_6409 ();
 sky130_fd_sc_hd__decap_3 PHY_6410 ();
 sky130_fd_sc_hd__decap_3 PHY_6411 ();
 sky130_fd_sc_hd__decap_3 PHY_6412 ();
 sky130_fd_sc_hd__decap_3 PHY_6413 ();
 sky130_fd_sc_hd__decap_3 PHY_6414 ();
 sky130_fd_sc_hd__decap_3 PHY_6415 ();
 sky130_fd_sc_hd__decap_3 PHY_6416 ();
 sky130_fd_sc_hd__decap_3 PHY_6417 ();
 sky130_fd_sc_hd__decap_3 PHY_6418 ();
 sky130_fd_sc_hd__decap_3 PHY_6419 ();
 sky130_fd_sc_hd__decap_3 PHY_6420 ();
 sky130_fd_sc_hd__decap_3 PHY_6421 ();
 sky130_fd_sc_hd__decap_3 PHY_6422 ();
 sky130_fd_sc_hd__decap_3 PHY_6423 ();
 sky130_fd_sc_hd__decap_3 PHY_6424 ();
 sky130_fd_sc_hd__decap_3 PHY_6425 ();
 sky130_fd_sc_hd__decap_3 PHY_6426 ();
 sky130_fd_sc_hd__decap_3 PHY_6427 ();
 sky130_fd_sc_hd__decap_3 PHY_6428 ();
 sky130_fd_sc_hd__decap_3 PHY_6429 ();
 sky130_fd_sc_hd__decap_3 PHY_6430 ();
 sky130_fd_sc_hd__decap_3 PHY_6431 ();
 sky130_fd_sc_hd__decap_3 PHY_6432 ();
 sky130_fd_sc_hd__decap_3 PHY_6433 ();
 sky130_fd_sc_hd__decap_3 PHY_6434 ();
 sky130_fd_sc_hd__decap_3 PHY_6435 ();
 sky130_fd_sc_hd__decap_3 PHY_6436 ();
 sky130_fd_sc_hd__decap_3 PHY_6437 ();
 sky130_fd_sc_hd__decap_3 PHY_6438 ();
 sky130_fd_sc_hd__decap_3 PHY_6439 ();
 sky130_fd_sc_hd__decap_3 PHY_6440 ();
 sky130_fd_sc_hd__decap_3 PHY_6441 ();
 sky130_fd_sc_hd__decap_3 PHY_6442 ();
 sky130_fd_sc_hd__decap_3 PHY_6443 ();
 sky130_fd_sc_hd__decap_3 PHY_6444 ();
 sky130_fd_sc_hd__decap_3 PHY_6445 ();
 sky130_fd_sc_hd__decap_3 PHY_6446 ();
 sky130_fd_sc_hd__decap_3 PHY_6447 ();
 sky130_fd_sc_hd__decap_3 PHY_6448 ();
 sky130_fd_sc_hd__decap_3 PHY_6449 ();
 sky130_fd_sc_hd__decap_3 PHY_6450 ();
 sky130_fd_sc_hd__decap_3 PHY_6451 ();
 sky130_fd_sc_hd__decap_3 PHY_6452 ();
 sky130_fd_sc_hd__decap_3 PHY_6453 ();
 sky130_fd_sc_hd__decap_3 PHY_6454 ();
 sky130_fd_sc_hd__decap_3 PHY_6455 ();
 sky130_fd_sc_hd__decap_3 PHY_6456 ();
 sky130_fd_sc_hd__decap_3 PHY_6457 ();
 sky130_fd_sc_hd__decap_3 PHY_6458 ();
 sky130_fd_sc_hd__decap_3 PHY_6459 ();
 sky130_fd_sc_hd__decap_3 PHY_6460 ();
 sky130_fd_sc_hd__decap_3 PHY_6461 ();
 sky130_fd_sc_hd__decap_3 PHY_6462 ();
 sky130_fd_sc_hd__decap_3 PHY_6463 ();
 sky130_fd_sc_hd__decap_3 PHY_6464 ();
 sky130_fd_sc_hd__decap_3 PHY_6465 ();
 sky130_fd_sc_hd__decap_3 PHY_6466 ();
 sky130_fd_sc_hd__decap_3 PHY_6467 ();
 sky130_fd_sc_hd__decap_3 PHY_6468 ();
 sky130_fd_sc_hd__decap_3 PHY_6469 ();
 sky130_fd_sc_hd__decap_3 PHY_6470 ();
 sky130_fd_sc_hd__decap_3 PHY_6471 ();
 sky130_fd_sc_hd__decap_3 PHY_6472 ();
 sky130_fd_sc_hd__decap_3 PHY_6473 ();
 sky130_fd_sc_hd__decap_3 PHY_6474 ();
 sky130_fd_sc_hd__decap_3 PHY_6475 ();
 sky130_fd_sc_hd__decap_3 PHY_6476 ();
 sky130_fd_sc_hd__decap_3 PHY_6477 ();
 sky130_fd_sc_hd__decap_3 PHY_6478 ();
 sky130_fd_sc_hd__decap_3 PHY_6479 ();
 sky130_fd_sc_hd__decap_3 PHY_6480 ();
 sky130_fd_sc_hd__decap_3 PHY_6481 ();
 sky130_fd_sc_hd__decap_3 PHY_6482 ();
 sky130_fd_sc_hd__decap_3 PHY_6483 ();
 sky130_fd_sc_hd__decap_3 PHY_6484 ();
 sky130_fd_sc_hd__decap_3 PHY_6485 ();
 sky130_fd_sc_hd__decap_3 PHY_6486 ();
 sky130_fd_sc_hd__decap_3 PHY_6487 ();
 sky130_fd_sc_hd__decap_3 PHY_6488 ();
 sky130_fd_sc_hd__decap_3 PHY_6489 ();
 sky130_fd_sc_hd__decap_3 PHY_6490 ();
 sky130_fd_sc_hd__decap_3 PHY_6491 ();
 sky130_fd_sc_hd__decap_3 PHY_6492 ();
 sky130_fd_sc_hd__decap_3 PHY_6493 ();
 sky130_fd_sc_hd__decap_3 PHY_6494 ();
 sky130_fd_sc_hd__decap_3 PHY_6495 ();
 sky130_fd_sc_hd__decap_3 PHY_6496 ();
 sky130_fd_sc_hd__decap_3 PHY_6497 ();
 sky130_fd_sc_hd__decap_3 PHY_6498 ();
 sky130_fd_sc_hd__decap_3 PHY_6499 ();
 sky130_fd_sc_hd__decap_3 PHY_6500 ();
 sky130_fd_sc_hd__decap_3 PHY_6501 ();
 sky130_fd_sc_hd__decap_3 PHY_6502 ();
 sky130_fd_sc_hd__decap_3 PHY_6503 ();
 sky130_fd_sc_hd__decap_3 PHY_6504 ();
 sky130_fd_sc_hd__decap_3 PHY_6505 ();
 sky130_fd_sc_hd__decap_3 PHY_6506 ();
 sky130_fd_sc_hd__decap_3 PHY_6507 ();
 sky130_fd_sc_hd__decap_3 PHY_6508 ();
 sky130_fd_sc_hd__decap_3 PHY_6509 ();
 sky130_fd_sc_hd__decap_3 PHY_6510 ();
 sky130_fd_sc_hd__decap_3 PHY_6511 ();
 sky130_fd_sc_hd__decap_3 PHY_6512 ();
 sky130_fd_sc_hd__decap_3 PHY_6513 ();
 sky130_fd_sc_hd__decap_3 PHY_6514 ();
 sky130_fd_sc_hd__decap_3 PHY_6515 ();
 sky130_fd_sc_hd__decap_3 PHY_6516 ();
 sky130_fd_sc_hd__decap_3 PHY_6517 ();
 sky130_fd_sc_hd__decap_3 PHY_6518 ();
 sky130_fd_sc_hd__decap_3 PHY_6519 ();
 sky130_fd_sc_hd__decap_3 PHY_6520 ();
 sky130_fd_sc_hd__decap_3 PHY_6521 ();
 sky130_fd_sc_hd__decap_3 PHY_6522 ();
 sky130_fd_sc_hd__decap_3 PHY_6523 ();
 sky130_fd_sc_hd__decap_3 PHY_6524 ();
 sky130_fd_sc_hd__decap_3 PHY_6525 ();
 sky130_fd_sc_hd__decap_3 PHY_6526 ();
 sky130_fd_sc_hd__decap_3 PHY_6527 ();
 sky130_fd_sc_hd__decap_3 PHY_6528 ();
 sky130_fd_sc_hd__decap_3 PHY_6529 ();
 sky130_fd_sc_hd__decap_3 PHY_6530 ();
 sky130_fd_sc_hd__decap_3 PHY_6531 ();
 sky130_fd_sc_hd__decap_3 PHY_6532 ();
 sky130_fd_sc_hd__decap_3 PHY_6533 ();
 sky130_fd_sc_hd__decap_3 PHY_6534 ();
 sky130_fd_sc_hd__decap_3 PHY_6535 ();
 sky130_fd_sc_hd__decap_3 PHY_6536 ();
 sky130_fd_sc_hd__decap_3 PHY_6537 ();
 sky130_fd_sc_hd__decap_3 PHY_6538 ();
 sky130_fd_sc_hd__decap_3 PHY_6539 ();
 sky130_fd_sc_hd__decap_3 PHY_6540 ();
 sky130_fd_sc_hd__decap_3 PHY_6541 ();
 sky130_fd_sc_hd__decap_3 PHY_6542 ();
 sky130_fd_sc_hd__decap_3 PHY_6543 ();
 sky130_fd_sc_hd__decap_3 PHY_6544 ();
 sky130_fd_sc_hd__decap_3 PHY_6545 ();
 sky130_fd_sc_hd__decap_3 PHY_6546 ();
 sky130_fd_sc_hd__decap_3 PHY_6547 ();
 sky130_fd_sc_hd__decap_3 PHY_6548 ();
 sky130_fd_sc_hd__decap_3 PHY_6549 ();
 sky130_fd_sc_hd__decap_3 PHY_6550 ();
 sky130_fd_sc_hd__decap_3 PHY_6551 ();
 sky130_fd_sc_hd__decap_3 PHY_6552 ();
 sky130_fd_sc_hd__decap_3 PHY_6553 ();
 sky130_fd_sc_hd__decap_3 PHY_6554 ();
 sky130_fd_sc_hd__decap_3 PHY_6555 ();
 sky130_fd_sc_hd__decap_3 PHY_6556 ();
 sky130_fd_sc_hd__decap_3 PHY_6557 ();
 sky130_fd_sc_hd__decap_3 PHY_6558 ();
 sky130_fd_sc_hd__decap_3 PHY_6559 ();
 sky130_fd_sc_hd__decap_3 PHY_6560 ();
 sky130_fd_sc_hd__decap_3 PHY_6561 ();
 sky130_fd_sc_hd__decap_3 PHY_6562 ();
 sky130_fd_sc_hd__decap_3 PHY_6563 ();
 sky130_fd_sc_hd__decap_3 PHY_6564 ();
 sky130_fd_sc_hd__decap_3 PHY_6565 ();
 sky130_fd_sc_hd__decap_3 PHY_6566 ();
 sky130_fd_sc_hd__decap_3 PHY_6567 ();
 sky130_fd_sc_hd__decap_3 PHY_6568 ();
 sky130_fd_sc_hd__decap_3 PHY_6569 ();
 sky130_fd_sc_hd__decap_3 PHY_6570 ();
 sky130_fd_sc_hd__decap_3 PHY_6571 ();
 sky130_fd_sc_hd__decap_3 PHY_6572 ();
 sky130_fd_sc_hd__decap_3 PHY_6573 ();
 sky130_fd_sc_hd__decap_3 PHY_6574 ();
 sky130_fd_sc_hd__decap_3 PHY_6575 ();
 sky130_fd_sc_hd__decap_3 PHY_6576 ();
 sky130_fd_sc_hd__decap_3 PHY_6577 ();
 sky130_fd_sc_hd__decap_3 PHY_6578 ();
 sky130_fd_sc_hd__decap_3 PHY_6579 ();
 sky130_fd_sc_hd__decap_3 PHY_6580 ();
 sky130_fd_sc_hd__decap_3 PHY_6581 ();
 sky130_fd_sc_hd__decap_3 PHY_6582 ();
 sky130_fd_sc_hd__decap_3 PHY_6583 ();
 sky130_fd_sc_hd__decap_3 PHY_6584 ();
 sky130_fd_sc_hd__decap_3 PHY_6585 ();
 sky130_fd_sc_hd__decap_3 PHY_6586 ();
 sky130_fd_sc_hd__decap_3 PHY_6587 ();
 sky130_fd_sc_hd__decap_3 PHY_6588 ();
 sky130_fd_sc_hd__decap_3 PHY_6589 ();
 sky130_fd_sc_hd__decap_3 PHY_6590 ();
 sky130_fd_sc_hd__decap_3 PHY_6591 ();
 sky130_fd_sc_hd__decap_3 PHY_6592 ();
 sky130_fd_sc_hd__decap_3 PHY_6593 ();
 sky130_fd_sc_hd__decap_3 PHY_6594 ();
 sky130_fd_sc_hd__decap_3 PHY_6595 ();
 sky130_fd_sc_hd__decap_3 PHY_6596 ();
 sky130_fd_sc_hd__decap_3 PHY_6597 ();
 sky130_fd_sc_hd__decap_3 PHY_6598 ();
 sky130_fd_sc_hd__decap_3 PHY_6599 ();
 sky130_fd_sc_hd__decap_3 PHY_6600 ();
 sky130_fd_sc_hd__decap_3 PHY_6601 ();
 sky130_fd_sc_hd__decap_3 PHY_6602 ();
 sky130_fd_sc_hd__decap_3 PHY_6603 ();
 sky130_fd_sc_hd__decap_3 PHY_6604 ();
 sky130_fd_sc_hd__decap_3 PHY_6605 ();
 sky130_fd_sc_hd__decap_3 PHY_6606 ();
 sky130_fd_sc_hd__decap_3 PHY_6607 ();
 sky130_fd_sc_hd__decap_3 PHY_6608 ();
 sky130_fd_sc_hd__decap_3 PHY_6609 ();
 sky130_fd_sc_hd__decap_3 PHY_6610 ();
 sky130_fd_sc_hd__decap_3 PHY_6611 ();
 sky130_fd_sc_hd__decap_3 PHY_6612 ();
 sky130_fd_sc_hd__decap_3 PHY_6613 ();
 sky130_fd_sc_hd__decap_3 PHY_6614 ();
 sky130_fd_sc_hd__decap_3 PHY_6615 ();
 sky130_fd_sc_hd__decap_3 PHY_6616 ();
 sky130_fd_sc_hd__decap_3 PHY_6617 ();
 sky130_fd_sc_hd__decap_3 PHY_6618 ();
 sky130_fd_sc_hd__decap_3 PHY_6619 ();
 sky130_fd_sc_hd__decap_3 PHY_6620 ();
 sky130_fd_sc_hd__decap_3 PHY_6621 ();
 sky130_fd_sc_hd__decap_3 PHY_6622 ();
 sky130_fd_sc_hd__decap_3 PHY_6623 ();
 sky130_fd_sc_hd__decap_3 PHY_6624 ();
 sky130_fd_sc_hd__decap_3 PHY_6625 ();
 sky130_fd_sc_hd__decap_3 PHY_6626 ();
 sky130_fd_sc_hd__decap_3 PHY_6627 ();
 sky130_fd_sc_hd__decap_3 PHY_6628 ();
 sky130_fd_sc_hd__decap_3 PHY_6629 ();
 sky130_fd_sc_hd__decap_3 PHY_6630 ();
 sky130_fd_sc_hd__decap_3 PHY_6631 ();
 sky130_fd_sc_hd__decap_3 PHY_6632 ();
 sky130_fd_sc_hd__decap_3 PHY_6633 ();
 sky130_fd_sc_hd__decap_3 PHY_6634 ();
 sky130_fd_sc_hd__decap_3 PHY_6635 ();
 sky130_fd_sc_hd__decap_3 PHY_6636 ();
 sky130_fd_sc_hd__decap_3 PHY_6637 ();
 sky130_fd_sc_hd__decap_3 PHY_6638 ();
 sky130_fd_sc_hd__decap_3 PHY_6639 ();
 sky130_fd_sc_hd__decap_3 PHY_6640 ();
 sky130_fd_sc_hd__decap_3 PHY_6641 ();
 sky130_fd_sc_hd__decap_3 PHY_6642 ();
 sky130_fd_sc_hd__decap_3 PHY_6643 ();
 sky130_fd_sc_hd__decap_3 PHY_6644 ();
 sky130_fd_sc_hd__decap_3 PHY_6645 ();
 sky130_fd_sc_hd__decap_3 PHY_6646 ();
 sky130_fd_sc_hd__decap_3 PHY_6647 ();
 sky130_fd_sc_hd__decap_3 PHY_6648 ();
 sky130_fd_sc_hd__decap_3 PHY_6649 ();
 sky130_fd_sc_hd__decap_3 PHY_6650 ();
 sky130_fd_sc_hd__decap_3 PHY_6651 ();
 sky130_fd_sc_hd__decap_3 PHY_6652 ();
 sky130_fd_sc_hd__decap_3 PHY_6653 ();
 sky130_fd_sc_hd__decap_3 PHY_6654 ();
 sky130_fd_sc_hd__decap_3 PHY_6655 ();
 sky130_fd_sc_hd__decap_3 PHY_6656 ();
 sky130_fd_sc_hd__decap_3 PHY_6657 ();
 sky130_fd_sc_hd__decap_3 PHY_6658 ();
 sky130_fd_sc_hd__decap_3 PHY_6659 ();
 sky130_fd_sc_hd__decap_3 PHY_6660 ();
 sky130_fd_sc_hd__decap_3 PHY_6661 ();
 sky130_fd_sc_hd__decap_3 PHY_6662 ();
 sky130_fd_sc_hd__decap_3 PHY_6663 ();
 sky130_fd_sc_hd__decap_3 PHY_6664 ();
 sky130_fd_sc_hd__decap_3 PHY_6665 ();
 sky130_fd_sc_hd__decap_3 PHY_6666 ();
 sky130_fd_sc_hd__decap_3 PHY_6667 ();
 sky130_fd_sc_hd__decap_3 PHY_6668 ();
 sky130_fd_sc_hd__decap_3 PHY_6669 ();
 sky130_fd_sc_hd__decap_3 PHY_6670 ();
 sky130_fd_sc_hd__decap_3 PHY_6671 ();
 sky130_fd_sc_hd__decap_3 PHY_6672 ();
 sky130_fd_sc_hd__decap_3 PHY_6673 ();
 sky130_fd_sc_hd__decap_3 PHY_6674 ();
 sky130_fd_sc_hd__decap_3 PHY_6675 ();
 sky130_fd_sc_hd__decap_3 PHY_6676 ();
 sky130_fd_sc_hd__decap_3 PHY_6677 ();
 sky130_fd_sc_hd__decap_3 PHY_6678 ();
 sky130_fd_sc_hd__decap_3 PHY_6679 ();
 sky130_fd_sc_hd__decap_3 PHY_6680 ();
 sky130_fd_sc_hd__decap_3 PHY_6681 ();
 sky130_fd_sc_hd__decap_3 PHY_6682 ();
 sky130_fd_sc_hd__decap_3 PHY_6683 ();
 sky130_fd_sc_hd__decap_3 PHY_6684 ();
 sky130_fd_sc_hd__decap_3 PHY_6685 ();
 sky130_fd_sc_hd__decap_3 PHY_6686 ();
 sky130_fd_sc_hd__decap_3 PHY_6687 ();
 sky130_fd_sc_hd__decap_3 PHY_6688 ();
 sky130_fd_sc_hd__decap_3 PHY_6689 ();
 sky130_fd_sc_hd__decap_3 PHY_6690 ();
 sky130_fd_sc_hd__decap_3 PHY_6691 ();
 sky130_fd_sc_hd__decap_3 PHY_6692 ();
 sky130_fd_sc_hd__decap_3 PHY_6693 ();
 sky130_fd_sc_hd__decap_3 PHY_6694 ();
 sky130_fd_sc_hd__decap_3 PHY_6695 ();
 sky130_fd_sc_hd__decap_3 PHY_6696 ();
 sky130_fd_sc_hd__decap_3 PHY_6697 ();
 sky130_fd_sc_hd__decap_3 PHY_6698 ();
 sky130_fd_sc_hd__decap_3 PHY_6699 ();
 sky130_fd_sc_hd__decap_3 PHY_6700 ();
 sky130_fd_sc_hd__decap_3 PHY_6701 ();
 sky130_fd_sc_hd__decap_3 PHY_6702 ();
 sky130_fd_sc_hd__decap_3 PHY_6703 ();
 sky130_fd_sc_hd__decap_3 PHY_6704 ();
 sky130_fd_sc_hd__decap_3 PHY_6705 ();
 sky130_fd_sc_hd__decap_3 PHY_6706 ();
 sky130_fd_sc_hd__decap_3 PHY_6707 ();
 sky130_fd_sc_hd__decap_3 PHY_6708 ();
 sky130_fd_sc_hd__decap_3 PHY_6709 ();
 sky130_fd_sc_hd__decap_3 PHY_6710 ();
 sky130_fd_sc_hd__decap_3 PHY_6711 ();
 sky130_fd_sc_hd__decap_3 PHY_6712 ();
 sky130_fd_sc_hd__decap_3 PHY_6713 ();
 sky130_fd_sc_hd__decap_3 PHY_6714 ();
 sky130_fd_sc_hd__decap_3 PHY_6715 ();
 sky130_fd_sc_hd__decap_3 PHY_6716 ();
 sky130_fd_sc_hd__decap_3 PHY_6717 ();
 sky130_fd_sc_hd__decap_3 PHY_6718 ();
 sky130_fd_sc_hd__decap_3 PHY_6719 ();
 sky130_fd_sc_hd__decap_3 PHY_6720 ();
 sky130_fd_sc_hd__decap_3 PHY_6721 ();
 sky130_fd_sc_hd__decap_3 PHY_6722 ();
 sky130_fd_sc_hd__decap_3 PHY_6723 ();
 sky130_fd_sc_hd__decap_3 PHY_6724 ();
 sky130_fd_sc_hd__decap_3 PHY_6725 ();
 sky130_fd_sc_hd__decap_3 PHY_6726 ();
 sky130_fd_sc_hd__decap_3 PHY_6727 ();
 sky130_fd_sc_hd__decap_3 PHY_6728 ();
 sky130_fd_sc_hd__decap_3 PHY_6729 ();
 sky130_fd_sc_hd__decap_3 PHY_6730 ();
 sky130_fd_sc_hd__decap_3 PHY_6731 ();
 sky130_fd_sc_hd__decap_3 PHY_6732 ();
 sky130_fd_sc_hd__decap_3 PHY_6733 ();
 sky130_fd_sc_hd__decap_3 PHY_6734 ();
 sky130_fd_sc_hd__decap_3 PHY_6735 ();
 sky130_fd_sc_hd__decap_3 PHY_6736 ();
 sky130_fd_sc_hd__decap_3 PHY_6737 ();
 sky130_fd_sc_hd__decap_3 PHY_6738 ();
 sky130_fd_sc_hd__decap_3 PHY_6739 ();
 sky130_fd_sc_hd__decap_3 PHY_6740 ();
 sky130_fd_sc_hd__decap_3 PHY_6741 ();
 sky130_fd_sc_hd__decap_3 PHY_6742 ();
 sky130_fd_sc_hd__decap_3 PHY_6743 ();
 sky130_fd_sc_hd__decap_3 PHY_6744 ();
 sky130_fd_sc_hd__decap_3 PHY_6745 ();
 sky130_fd_sc_hd__decap_3 PHY_6746 ();
 sky130_fd_sc_hd__decap_3 PHY_6747 ();
 sky130_fd_sc_hd__decap_3 PHY_6748 ();
 sky130_fd_sc_hd__decap_3 PHY_6749 ();
 sky130_fd_sc_hd__decap_3 PHY_6750 ();
 sky130_fd_sc_hd__decap_3 PHY_6751 ();
 sky130_fd_sc_hd__decap_3 PHY_6752 ();
 sky130_fd_sc_hd__decap_3 PHY_6753 ();
 sky130_fd_sc_hd__decap_3 PHY_6754 ();
 sky130_fd_sc_hd__decap_3 PHY_6755 ();
 sky130_fd_sc_hd__decap_3 PHY_6756 ();
 sky130_fd_sc_hd__decap_3 PHY_6757 ();
 sky130_fd_sc_hd__decap_3 PHY_6758 ();
 sky130_fd_sc_hd__decap_3 PHY_6759 ();
 sky130_fd_sc_hd__decap_3 PHY_6760 ();
 sky130_fd_sc_hd__decap_3 PHY_6761 ();
 sky130_fd_sc_hd__decap_3 PHY_6762 ();
 sky130_fd_sc_hd__decap_3 PHY_6763 ();
 sky130_fd_sc_hd__decap_3 PHY_6764 ();
 sky130_fd_sc_hd__decap_3 PHY_6765 ();
 sky130_fd_sc_hd__decap_3 PHY_6766 ();
 sky130_fd_sc_hd__decap_3 PHY_6767 ();
 sky130_fd_sc_hd__decap_3 PHY_6768 ();
 sky130_fd_sc_hd__decap_3 PHY_6769 ();
 sky130_fd_sc_hd__decap_3 PHY_6770 ();
 sky130_fd_sc_hd__decap_3 PHY_6771 ();
 sky130_fd_sc_hd__decap_3 PHY_6772 ();
 sky130_fd_sc_hd__decap_3 PHY_6773 ();
 sky130_fd_sc_hd__decap_3 PHY_6774 ();
 sky130_fd_sc_hd__decap_3 PHY_6775 ();
 sky130_fd_sc_hd__decap_3 PHY_6776 ();
 sky130_fd_sc_hd__decap_3 PHY_6777 ();
 sky130_fd_sc_hd__decap_3 PHY_6778 ();
 sky130_fd_sc_hd__decap_3 PHY_6779 ();
 sky130_fd_sc_hd__decap_3 PHY_6780 ();
 sky130_fd_sc_hd__decap_3 PHY_6781 ();
 sky130_fd_sc_hd__decap_3 PHY_6782 ();
 sky130_fd_sc_hd__decap_3 PHY_6783 ();
 sky130_fd_sc_hd__decap_3 PHY_6784 ();
 sky130_fd_sc_hd__decap_3 PHY_6785 ();
 sky130_fd_sc_hd__decap_3 PHY_6786 ();
 sky130_fd_sc_hd__decap_3 PHY_6787 ();
 sky130_fd_sc_hd__decap_3 PHY_6788 ();
 sky130_fd_sc_hd__decap_3 PHY_6789 ();
 sky130_fd_sc_hd__decap_3 PHY_6790 ();
 sky130_fd_sc_hd__decap_3 PHY_6791 ();
 sky130_fd_sc_hd__decap_3 PHY_6792 ();
 sky130_fd_sc_hd__decap_3 PHY_6793 ();
 sky130_fd_sc_hd__decap_3 PHY_6794 ();
 sky130_fd_sc_hd__decap_3 PHY_6795 ();
 sky130_fd_sc_hd__decap_3 PHY_6796 ();
 sky130_fd_sc_hd__decap_3 PHY_6797 ();
 sky130_fd_sc_hd__decap_3 PHY_6798 ();
 sky130_fd_sc_hd__decap_3 PHY_6799 ();
 sky130_fd_sc_hd__decap_3 PHY_6800 ();
 sky130_fd_sc_hd__decap_3 PHY_6801 ();
 sky130_fd_sc_hd__decap_3 PHY_6802 ();
 sky130_fd_sc_hd__decap_3 PHY_6803 ();
 sky130_fd_sc_hd__decap_3 PHY_6804 ();
 sky130_fd_sc_hd__decap_3 PHY_6805 ();
 sky130_fd_sc_hd__decap_3 PHY_6806 ();
 sky130_fd_sc_hd__decap_3 PHY_6807 ();
 sky130_fd_sc_hd__decap_3 PHY_6808 ();
 sky130_fd_sc_hd__decap_3 PHY_6809 ();
 sky130_fd_sc_hd__decap_3 PHY_6810 ();
 sky130_fd_sc_hd__decap_3 PHY_6811 ();
 sky130_fd_sc_hd__decap_3 PHY_6812 ();
 sky130_fd_sc_hd__decap_3 PHY_6813 ();
 sky130_fd_sc_hd__decap_3 PHY_6814 ();
 sky130_fd_sc_hd__decap_3 PHY_6815 ();
 sky130_fd_sc_hd__decap_3 PHY_6816 ();
 sky130_fd_sc_hd__decap_3 PHY_6817 ();
 sky130_fd_sc_hd__decap_3 PHY_6818 ();
 sky130_fd_sc_hd__decap_3 PHY_6819 ();
 sky130_fd_sc_hd__decap_3 PHY_6820 ();
 sky130_fd_sc_hd__decap_3 PHY_6821 ();
 sky130_fd_sc_hd__decap_3 PHY_6822 ();
 sky130_fd_sc_hd__decap_3 PHY_6823 ();
 sky130_fd_sc_hd__decap_3 PHY_6824 ();
 sky130_fd_sc_hd__decap_3 PHY_6825 ();
 sky130_fd_sc_hd__decap_3 PHY_6826 ();
 sky130_fd_sc_hd__decap_3 PHY_6827 ();
 sky130_fd_sc_hd__decap_3 PHY_6828 ();
 sky130_fd_sc_hd__decap_3 PHY_6829 ();
 sky130_fd_sc_hd__decap_3 PHY_6830 ();
 sky130_fd_sc_hd__decap_3 PHY_6831 ();
 sky130_fd_sc_hd__decap_3 PHY_6832 ();
 sky130_fd_sc_hd__decap_3 PHY_6833 ();
 sky130_fd_sc_hd__decap_3 PHY_6834 ();
 sky130_fd_sc_hd__decap_3 PHY_6835 ();
 sky130_fd_sc_hd__decap_3 PHY_6836 ();
 sky130_fd_sc_hd__decap_3 PHY_6837 ();
 sky130_fd_sc_hd__decap_3 PHY_6838 ();
 sky130_fd_sc_hd__decap_3 PHY_6839 ();
 sky130_fd_sc_hd__decap_3 PHY_6840 ();
 sky130_fd_sc_hd__decap_3 PHY_6841 ();
 sky130_fd_sc_hd__decap_3 PHY_6842 ();
 sky130_fd_sc_hd__decap_3 PHY_6843 ();
 sky130_fd_sc_hd__decap_3 PHY_6844 ();
 sky130_fd_sc_hd__decap_3 PHY_6845 ();
 sky130_fd_sc_hd__decap_3 PHY_6846 ();
 sky130_fd_sc_hd__decap_3 PHY_6847 ();
 sky130_fd_sc_hd__decap_3 PHY_6848 ();
 sky130_fd_sc_hd__decap_3 PHY_6849 ();
 sky130_fd_sc_hd__decap_3 PHY_6850 ();
 sky130_fd_sc_hd__decap_3 PHY_6851 ();
 sky130_fd_sc_hd__decap_3 PHY_6852 ();
 sky130_fd_sc_hd__decap_3 PHY_6853 ();
 sky130_fd_sc_hd__decap_3 PHY_6854 ();
 sky130_fd_sc_hd__decap_3 PHY_6855 ();
 sky130_fd_sc_hd__decap_3 PHY_6856 ();
 sky130_fd_sc_hd__decap_3 PHY_6857 ();
 sky130_fd_sc_hd__decap_3 PHY_6858 ();
 sky130_fd_sc_hd__decap_3 PHY_6859 ();
 sky130_fd_sc_hd__decap_3 PHY_6860 ();
 sky130_fd_sc_hd__decap_3 PHY_6861 ();
 sky130_fd_sc_hd__decap_3 PHY_6862 ();
 sky130_fd_sc_hd__decap_3 PHY_6863 ();
 sky130_fd_sc_hd__decap_3 PHY_6864 ();
 sky130_fd_sc_hd__decap_3 PHY_6865 ();
 sky130_fd_sc_hd__decap_3 PHY_6866 ();
 sky130_fd_sc_hd__decap_3 PHY_6867 ();
 sky130_fd_sc_hd__decap_3 PHY_6868 ();
 sky130_fd_sc_hd__decap_3 PHY_6869 ();
 sky130_fd_sc_hd__decap_3 PHY_6870 ();
 sky130_fd_sc_hd__decap_3 PHY_6871 ();
 sky130_fd_sc_hd__decap_3 PHY_6872 ();
 sky130_fd_sc_hd__decap_3 PHY_6873 ();
 sky130_fd_sc_hd__decap_3 PHY_6874 ();
 sky130_fd_sc_hd__decap_3 PHY_6875 ();
 sky130_fd_sc_hd__decap_3 PHY_6876 ();
 sky130_fd_sc_hd__decap_3 PHY_6877 ();
 sky130_fd_sc_hd__decap_3 PHY_6878 ();
 sky130_fd_sc_hd__decap_3 PHY_6879 ();
 sky130_fd_sc_hd__decap_3 PHY_6880 ();
 sky130_fd_sc_hd__decap_3 PHY_6881 ();
 sky130_fd_sc_hd__decap_3 PHY_6882 ();
 sky130_fd_sc_hd__decap_3 PHY_6883 ();
 sky130_fd_sc_hd__decap_3 PHY_6884 ();
 sky130_fd_sc_hd__decap_3 PHY_6885 ();
 sky130_fd_sc_hd__decap_3 PHY_6886 ();
 sky130_fd_sc_hd__decap_3 PHY_6887 ();
 sky130_fd_sc_hd__decap_3 PHY_6888 ();
 sky130_fd_sc_hd__decap_3 PHY_6889 ();
 sky130_fd_sc_hd__decap_3 PHY_6890 ();
 sky130_fd_sc_hd__decap_3 PHY_6891 ();
 sky130_fd_sc_hd__decap_3 PHY_6892 ();
 sky130_fd_sc_hd__decap_3 PHY_6893 ();
 sky130_fd_sc_hd__decap_3 PHY_6894 ();
 sky130_fd_sc_hd__decap_3 PHY_6895 ();
 sky130_fd_sc_hd__decap_3 PHY_6896 ();
 sky130_fd_sc_hd__decap_3 PHY_6897 ();
 sky130_fd_sc_hd__decap_3 PHY_6898 ();
 sky130_fd_sc_hd__decap_3 PHY_6899 ();
 sky130_fd_sc_hd__decap_3 PHY_6900 ();
 sky130_fd_sc_hd__decap_3 PHY_6901 ();
 sky130_fd_sc_hd__decap_3 PHY_6902 ();
 sky130_fd_sc_hd__decap_3 PHY_6903 ();
 sky130_fd_sc_hd__decap_3 PHY_6904 ();
 sky130_fd_sc_hd__decap_3 PHY_6905 ();
 sky130_fd_sc_hd__decap_3 PHY_6906 ();
 sky130_fd_sc_hd__decap_3 PHY_6907 ();
 sky130_fd_sc_hd__decap_3 PHY_6908 ();
 sky130_fd_sc_hd__decap_3 PHY_6909 ();
 sky130_fd_sc_hd__decap_3 PHY_6910 ();
 sky130_fd_sc_hd__decap_3 PHY_6911 ();
 sky130_fd_sc_hd__decap_3 PHY_6912 ();
 sky130_fd_sc_hd__decap_3 PHY_6913 ();
 sky130_fd_sc_hd__decap_3 PHY_6914 ();
 sky130_fd_sc_hd__decap_3 PHY_6915 ();
 sky130_fd_sc_hd__decap_3 PHY_6916 ();
 sky130_fd_sc_hd__decap_3 PHY_6917 ();
 sky130_fd_sc_hd__decap_3 PHY_6918 ();
 sky130_fd_sc_hd__decap_3 PHY_6919 ();
 sky130_fd_sc_hd__decap_3 PHY_6920 ();
 sky130_fd_sc_hd__decap_3 PHY_6921 ();
 sky130_fd_sc_hd__decap_3 PHY_6922 ();
 sky130_fd_sc_hd__decap_3 PHY_6923 ();
 sky130_fd_sc_hd__decap_3 PHY_6924 ();
 sky130_fd_sc_hd__decap_3 PHY_6925 ();
 sky130_fd_sc_hd__decap_3 PHY_6926 ();
 sky130_fd_sc_hd__decap_3 PHY_6927 ();
 sky130_fd_sc_hd__decap_3 PHY_6928 ();
 sky130_fd_sc_hd__decap_3 PHY_6929 ();
 sky130_fd_sc_hd__decap_3 PHY_6930 ();
 sky130_fd_sc_hd__decap_3 PHY_6931 ();
 sky130_fd_sc_hd__decap_3 PHY_6932 ();
 sky130_fd_sc_hd__decap_3 PHY_6933 ();
 sky130_fd_sc_hd__decap_3 PHY_6934 ();
 sky130_fd_sc_hd__decap_3 PHY_6935 ();
 sky130_fd_sc_hd__decap_3 PHY_6936 ();
 sky130_fd_sc_hd__decap_3 PHY_6937 ();
 sky130_fd_sc_hd__decap_3 PHY_6938 ();
 sky130_fd_sc_hd__decap_3 PHY_6939 ();
 sky130_fd_sc_hd__decap_3 PHY_6940 ();
 sky130_fd_sc_hd__decap_3 PHY_6941 ();
 sky130_fd_sc_hd__decap_3 PHY_6942 ();
 sky130_fd_sc_hd__decap_3 PHY_6943 ();
 sky130_fd_sc_hd__decap_3 PHY_6944 ();
 sky130_fd_sc_hd__decap_3 PHY_6945 ();
 sky130_fd_sc_hd__decap_3 PHY_6946 ();
 sky130_fd_sc_hd__decap_3 PHY_6947 ();
 sky130_fd_sc_hd__decap_3 PHY_6948 ();
 sky130_fd_sc_hd__decap_3 PHY_6949 ();
 sky130_fd_sc_hd__decap_3 PHY_6950 ();
 sky130_fd_sc_hd__decap_3 PHY_6951 ();
 sky130_fd_sc_hd__decap_3 PHY_6952 ();
 sky130_fd_sc_hd__decap_3 PHY_6953 ();
 sky130_fd_sc_hd__decap_3 PHY_6954 ();
 sky130_fd_sc_hd__decap_3 PHY_6955 ();
 sky130_fd_sc_hd__decap_3 PHY_6956 ();
 sky130_fd_sc_hd__decap_3 PHY_6957 ();
 sky130_fd_sc_hd__decap_3 PHY_6958 ();
 sky130_fd_sc_hd__decap_3 PHY_6959 ();
 sky130_fd_sc_hd__decap_3 PHY_6960 ();
 sky130_fd_sc_hd__decap_3 PHY_6961 ();
 sky130_fd_sc_hd__decap_3 PHY_6962 ();
 sky130_fd_sc_hd__decap_3 PHY_6963 ();
 sky130_fd_sc_hd__decap_3 PHY_6964 ();
 sky130_fd_sc_hd__decap_3 PHY_6965 ();
 sky130_fd_sc_hd__decap_3 PHY_6966 ();
 sky130_fd_sc_hd__decap_3 PHY_6967 ();
 sky130_fd_sc_hd__decap_3 PHY_6968 ();
 sky130_fd_sc_hd__decap_3 PHY_6969 ();
 sky130_fd_sc_hd__decap_3 PHY_6970 ();
 sky130_fd_sc_hd__decap_3 PHY_6971 ();
 sky130_fd_sc_hd__decap_3 PHY_6972 ();
 sky130_fd_sc_hd__decap_3 PHY_6973 ();
 sky130_fd_sc_hd__decap_3 PHY_6974 ();
 sky130_fd_sc_hd__decap_3 PHY_6975 ();
 sky130_fd_sc_hd__decap_3 PHY_6976 ();
 sky130_fd_sc_hd__decap_3 PHY_6977 ();
 sky130_fd_sc_hd__decap_3 PHY_6978 ();
 sky130_fd_sc_hd__decap_3 PHY_6979 ();
 sky130_fd_sc_hd__decap_3 PHY_6980 ();
 sky130_fd_sc_hd__decap_3 PHY_6981 ();
 sky130_fd_sc_hd__decap_3 PHY_6982 ();
 sky130_fd_sc_hd__decap_3 PHY_6983 ();
 sky130_fd_sc_hd__decap_3 PHY_6984 ();
 sky130_fd_sc_hd__decap_3 PHY_6985 ();
 sky130_fd_sc_hd__decap_3 PHY_6986 ();
 sky130_fd_sc_hd__decap_3 PHY_6987 ();
 sky130_fd_sc_hd__decap_3 PHY_6988 ();
 sky130_fd_sc_hd__decap_3 PHY_6989 ();
 sky130_fd_sc_hd__decap_3 PHY_6990 ();
 sky130_fd_sc_hd__decap_3 PHY_6991 ();
 sky130_fd_sc_hd__decap_3 PHY_6992 ();
 sky130_fd_sc_hd__decap_3 PHY_6993 ();
 sky130_fd_sc_hd__decap_3 PHY_6994 ();
 sky130_fd_sc_hd__decap_3 PHY_6995 ();
 sky130_fd_sc_hd__decap_3 PHY_6996 ();
 sky130_fd_sc_hd__decap_3 PHY_6997 ();
 sky130_fd_sc_hd__decap_3 PHY_6998 ();
 sky130_fd_sc_hd__decap_3 PHY_6999 ();
 sky130_fd_sc_hd__decap_3 PHY_7000 ();
 sky130_fd_sc_hd__decap_3 PHY_7001 ();
 sky130_fd_sc_hd__decap_3 PHY_7002 ();
 sky130_fd_sc_hd__decap_3 PHY_7003 ();
 sky130_fd_sc_hd__decap_3 PHY_7004 ();
 sky130_fd_sc_hd__decap_3 PHY_7005 ();
 sky130_fd_sc_hd__decap_3 PHY_7006 ();
 sky130_fd_sc_hd__decap_3 PHY_7007 ();
 sky130_fd_sc_hd__decap_3 PHY_7008 ();
 sky130_fd_sc_hd__decap_3 PHY_7009 ();
 sky130_fd_sc_hd__decap_3 PHY_7010 ();
 sky130_fd_sc_hd__decap_3 PHY_7011 ();
 sky130_fd_sc_hd__decap_3 PHY_7012 ();
 sky130_fd_sc_hd__decap_3 PHY_7013 ();
 sky130_fd_sc_hd__decap_3 PHY_7014 ();
 sky130_fd_sc_hd__decap_3 PHY_7015 ();
 sky130_fd_sc_hd__decap_3 PHY_7016 ();
 sky130_fd_sc_hd__decap_3 PHY_7017 ();
 sky130_fd_sc_hd__decap_3 PHY_7018 ();
 sky130_fd_sc_hd__decap_3 PHY_7019 ();
 sky130_fd_sc_hd__decap_3 PHY_7020 ();
 sky130_fd_sc_hd__decap_3 PHY_7021 ();
 sky130_fd_sc_hd__decap_3 PHY_7022 ();
 sky130_fd_sc_hd__decap_3 PHY_7023 ();
 sky130_fd_sc_hd__decap_3 PHY_7024 ();
 sky130_fd_sc_hd__decap_3 PHY_7025 ();
 sky130_fd_sc_hd__decap_3 PHY_7026 ();
 sky130_fd_sc_hd__decap_3 PHY_7027 ();
 sky130_fd_sc_hd__decap_3 PHY_7028 ();
 sky130_fd_sc_hd__decap_3 PHY_7029 ();
 sky130_fd_sc_hd__decap_3 PHY_7030 ();
 sky130_fd_sc_hd__decap_3 PHY_7031 ();
 sky130_fd_sc_hd__decap_3 PHY_7032 ();
 sky130_fd_sc_hd__decap_3 PHY_7033 ();
 sky130_fd_sc_hd__decap_3 PHY_7034 ();
 sky130_fd_sc_hd__decap_3 PHY_7035 ();
 sky130_fd_sc_hd__decap_3 PHY_7036 ();
 sky130_fd_sc_hd__decap_3 PHY_7037 ();
 sky130_fd_sc_hd__decap_3 PHY_7038 ();
 sky130_fd_sc_hd__decap_3 PHY_7039 ();
 sky130_fd_sc_hd__decap_3 PHY_7040 ();
 sky130_fd_sc_hd__decap_3 PHY_7041 ();
 sky130_fd_sc_hd__decap_3 PHY_7042 ();
 sky130_fd_sc_hd__decap_3 PHY_7043 ();
 sky130_fd_sc_hd__decap_3 PHY_7044 ();
 sky130_fd_sc_hd__decap_3 PHY_7045 ();
 sky130_fd_sc_hd__decap_3 PHY_7046 ();
 sky130_fd_sc_hd__decap_3 PHY_7047 ();
 sky130_fd_sc_hd__decap_3 PHY_7048 ();
 sky130_fd_sc_hd__decap_3 PHY_7049 ();
 sky130_fd_sc_hd__decap_3 PHY_7050 ();
 sky130_fd_sc_hd__decap_3 PHY_7051 ();
 sky130_fd_sc_hd__decap_3 PHY_7052 ();
 sky130_fd_sc_hd__decap_3 PHY_7053 ();
 sky130_fd_sc_hd__decap_3 PHY_7054 ();
 sky130_fd_sc_hd__decap_3 PHY_7055 ();
 sky130_fd_sc_hd__decap_3 PHY_7056 ();
 sky130_fd_sc_hd__decap_3 PHY_7057 ();
 sky130_fd_sc_hd__decap_3 PHY_7058 ();
 sky130_fd_sc_hd__decap_3 PHY_7059 ();
 sky130_fd_sc_hd__decap_3 PHY_7060 ();
 sky130_fd_sc_hd__decap_3 PHY_7061 ();
 sky130_fd_sc_hd__decap_3 PHY_7062 ();
 sky130_fd_sc_hd__decap_3 PHY_7063 ();
 sky130_fd_sc_hd__decap_3 PHY_7064 ();
 sky130_fd_sc_hd__decap_3 PHY_7065 ();
 sky130_fd_sc_hd__decap_3 PHY_7066 ();
 sky130_fd_sc_hd__decap_3 PHY_7067 ();
 sky130_fd_sc_hd__decap_3 PHY_7068 ();
 sky130_fd_sc_hd__decap_3 PHY_7069 ();
 sky130_fd_sc_hd__decap_3 PHY_7070 ();
 sky130_fd_sc_hd__decap_3 PHY_7071 ();
 sky130_fd_sc_hd__decap_3 PHY_7072 ();
 sky130_fd_sc_hd__decap_3 PHY_7073 ();
 sky130_fd_sc_hd__decap_3 PHY_7074 ();
 sky130_fd_sc_hd__decap_3 PHY_7075 ();
 sky130_fd_sc_hd__decap_3 PHY_7076 ();
 sky130_fd_sc_hd__decap_3 PHY_7077 ();
 sky130_fd_sc_hd__decap_3 PHY_7078 ();
 sky130_fd_sc_hd__decap_3 PHY_7079 ();
 sky130_fd_sc_hd__decap_3 PHY_7080 ();
 sky130_fd_sc_hd__decap_3 PHY_7081 ();
 sky130_fd_sc_hd__decap_3 PHY_7082 ();
 sky130_fd_sc_hd__decap_3 PHY_7083 ();
 sky130_fd_sc_hd__decap_3 PHY_7084 ();
 sky130_fd_sc_hd__decap_3 PHY_7085 ();
 sky130_fd_sc_hd__decap_3 PHY_7086 ();
 sky130_fd_sc_hd__decap_3 PHY_7087 ();
 sky130_fd_sc_hd__decap_3 PHY_7088 ();
 sky130_fd_sc_hd__decap_3 PHY_7089 ();
 sky130_fd_sc_hd__decap_3 PHY_7090 ();
 sky130_fd_sc_hd__decap_3 PHY_7091 ();
 sky130_fd_sc_hd__decap_3 PHY_7092 ();
 sky130_fd_sc_hd__decap_3 PHY_7093 ();
 sky130_fd_sc_hd__decap_3 PHY_7094 ();
 sky130_fd_sc_hd__decap_3 PHY_7095 ();
 sky130_fd_sc_hd__decap_3 PHY_7096 ();
 sky130_fd_sc_hd__decap_3 PHY_7097 ();
 sky130_fd_sc_hd__decap_3 PHY_7098 ();
 sky130_fd_sc_hd__decap_3 PHY_7099 ();
 sky130_fd_sc_hd__decap_3 PHY_7100 ();
 sky130_fd_sc_hd__decap_3 PHY_7101 ();
 sky130_fd_sc_hd__decap_3 PHY_7102 ();
 sky130_fd_sc_hd__decap_3 PHY_7103 ();
 sky130_fd_sc_hd__decap_3 PHY_7104 ();
 sky130_fd_sc_hd__decap_3 PHY_7105 ();
 sky130_fd_sc_hd__decap_3 PHY_7106 ();
 sky130_fd_sc_hd__decap_3 PHY_7107 ();
 sky130_fd_sc_hd__decap_3 PHY_7108 ();
 sky130_fd_sc_hd__decap_3 PHY_7109 ();
 sky130_fd_sc_hd__decap_3 PHY_7110 ();
 sky130_fd_sc_hd__decap_3 PHY_7111 ();
 sky130_fd_sc_hd__decap_3 PHY_7112 ();
 sky130_fd_sc_hd__decap_3 PHY_7113 ();
 sky130_fd_sc_hd__decap_3 PHY_7114 ();
 sky130_fd_sc_hd__decap_3 PHY_7115 ();
 sky130_fd_sc_hd__decap_3 PHY_7116 ();
 sky130_fd_sc_hd__decap_3 PHY_7117 ();
 sky130_fd_sc_hd__decap_3 PHY_7118 ();
 sky130_fd_sc_hd__decap_3 PHY_7119 ();
 sky130_fd_sc_hd__decap_3 PHY_7120 ();
 sky130_fd_sc_hd__decap_3 PHY_7121 ();
 sky130_fd_sc_hd__decap_3 PHY_7122 ();
 sky130_fd_sc_hd__decap_3 PHY_7123 ();
 sky130_fd_sc_hd__decap_3 PHY_7124 ();
 sky130_fd_sc_hd__decap_3 PHY_7125 ();
 sky130_fd_sc_hd__decap_3 PHY_7126 ();
 sky130_fd_sc_hd__decap_3 PHY_7127 ();
 sky130_fd_sc_hd__decap_3 PHY_7128 ();
 sky130_fd_sc_hd__decap_3 PHY_7129 ();
 sky130_fd_sc_hd__decap_3 PHY_7130 ();
 sky130_fd_sc_hd__decap_3 PHY_7131 ();
 sky130_fd_sc_hd__decap_3 PHY_7132 ();
 sky130_fd_sc_hd__decap_3 PHY_7133 ();
 sky130_fd_sc_hd__decap_3 PHY_7134 ();
 sky130_fd_sc_hd__decap_3 PHY_7135 ();
 sky130_fd_sc_hd__decap_3 PHY_7136 ();
 sky130_fd_sc_hd__decap_3 PHY_7137 ();
 sky130_fd_sc_hd__decap_3 PHY_7138 ();
 sky130_fd_sc_hd__decap_3 PHY_7139 ();
 sky130_fd_sc_hd__decap_3 PHY_7140 ();
 sky130_fd_sc_hd__decap_3 PHY_7141 ();
 sky130_fd_sc_hd__decap_3 PHY_7142 ();
 sky130_fd_sc_hd__decap_3 PHY_7143 ();
 sky130_fd_sc_hd__decap_3 PHY_7144 ();
 sky130_fd_sc_hd__decap_3 PHY_7145 ();
 sky130_fd_sc_hd__decap_3 PHY_7146 ();
 sky130_fd_sc_hd__decap_3 PHY_7147 ();
 sky130_fd_sc_hd__decap_3 PHY_7148 ();
 sky130_fd_sc_hd__decap_3 PHY_7149 ();
 sky130_fd_sc_hd__decap_3 PHY_7150 ();
 sky130_fd_sc_hd__decap_3 PHY_7151 ();
 sky130_fd_sc_hd__decap_3 PHY_7152 ();
 sky130_fd_sc_hd__decap_3 PHY_7153 ();
 sky130_fd_sc_hd__decap_3 PHY_7154 ();
 sky130_fd_sc_hd__decap_3 PHY_7155 ();
 sky130_fd_sc_hd__decap_3 PHY_7156 ();
 sky130_fd_sc_hd__decap_3 PHY_7157 ();
 sky130_fd_sc_hd__decap_3 PHY_7158 ();
 sky130_fd_sc_hd__decap_3 PHY_7159 ();
 sky130_fd_sc_hd__decap_3 PHY_7160 ();
 sky130_fd_sc_hd__decap_3 PHY_7161 ();
 sky130_fd_sc_hd__decap_3 PHY_7162 ();
 sky130_fd_sc_hd__decap_3 PHY_7163 ();
 sky130_fd_sc_hd__decap_3 PHY_7164 ();
 sky130_fd_sc_hd__decap_3 PHY_7165 ();
 sky130_fd_sc_hd__decap_3 PHY_7166 ();
 sky130_fd_sc_hd__decap_3 PHY_7167 ();
 sky130_fd_sc_hd__decap_3 PHY_7168 ();
 sky130_fd_sc_hd__decap_3 PHY_7169 ();
 sky130_fd_sc_hd__decap_3 PHY_7170 ();
 sky130_fd_sc_hd__decap_3 PHY_7171 ();
 sky130_fd_sc_hd__decap_3 PHY_7172 ();
 sky130_fd_sc_hd__decap_3 PHY_7173 ();
 sky130_fd_sc_hd__decap_3 PHY_7174 ();
 sky130_fd_sc_hd__decap_3 PHY_7175 ();
 sky130_fd_sc_hd__decap_3 PHY_7176 ();
 sky130_fd_sc_hd__decap_3 PHY_7177 ();
 sky130_fd_sc_hd__decap_3 PHY_7178 ();
 sky130_fd_sc_hd__decap_3 PHY_7179 ();
 sky130_fd_sc_hd__decap_3 PHY_7180 ();
 sky130_fd_sc_hd__decap_3 PHY_7181 ();
 sky130_fd_sc_hd__decap_3 PHY_7182 ();
 sky130_fd_sc_hd__decap_3 PHY_7183 ();
 sky130_fd_sc_hd__decap_3 PHY_7184 ();
 sky130_fd_sc_hd__decap_3 PHY_7185 ();
 sky130_fd_sc_hd__decap_3 PHY_7186 ();
 sky130_fd_sc_hd__decap_3 PHY_7187 ();
 sky130_fd_sc_hd__decap_3 PHY_7188 ();
 sky130_fd_sc_hd__decap_3 PHY_7189 ();
 sky130_fd_sc_hd__decap_3 PHY_7190 ();
 sky130_fd_sc_hd__decap_3 PHY_7191 ();
 sky130_fd_sc_hd__decap_3 PHY_7192 ();
 sky130_fd_sc_hd__decap_3 PHY_7193 ();
 sky130_fd_sc_hd__decap_3 PHY_7194 ();
 sky130_fd_sc_hd__decap_3 PHY_7195 ();
 sky130_fd_sc_hd__decap_3 PHY_7196 ();
 sky130_fd_sc_hd__decap_3 PHY_7197 ();
 sky130_fd_sc_hd__decap_3 PHY_7198 ();
 sky130_fd_sc_hd__decap_3 PHY_7199 ();
 sky130_fd_sc_hd__decap_3 PHY_7200 ();
 sky130_fd_sc_hd__decap_3 PHY_7201 ();
 sky130_fd_sc_hd__decap_3 PHY_7202 ();
 sky130_fd_sc_hd__decap_3 PHY_7203 ();
 sky130_fd_sc_hd__decap_3 PHY_7204 ();
 sky130_fd_sc_hd__decap_3 PHY_7205 ();
 sky130_fd_sc_hd__decap_3 PHY_7206 ();
 sky130_fd_sc_hd__decap_3 PHY_7207 ();
 sky130_fd_sc_hd__decap_3 PHY_7208 ();
 sky130_fd_sc_hd__decap_3 PHY_7209 ();
 sky130_fd_sc_hd__decap_3 PHY_7210 ();
 sky130_fd_sc_hd__decap_3 PHY_7211 ();
 sky130_fd_sc_hd__decap_3 PHY_7212 ();
 sky130_fd_sc_hd__decap_3 PHY_7213 ();
 sky130_fd_sc_hd__decap_3 PHY_7214 ();
 sky130_fd_sc_hd__decap_3 PHY_7215 ();
 sky130_fd_sc_hd__decap_3 PHY_7216 ();
 sky130_fd_sc_hd__decap_3 PHY_7217 ();
 sky130_fd_sc_hd__decap_3 PHY_7218 ();
 sky130_fd_sc_hd__decap_3 PHY_7219 ();
 sky130_fd_sc_hd__decap_3 PHY_7220 ();
 sky130_fd_sc_hd__decap_3 PHY_7221 ();
 sky130_fd_sc_hd__decap_3 PHY_7222 ();
 sky130_fd_sc_hd__decap_3 PHY_7223 ();
 sky130_fd_sc_hd__decap_3 PHY_7224 ();
 sky130_fd_sc_hd__decap_3 PHY_7225 ();
 sky130_fd_sc_hd__decap_3 PHY_7226 ();
 sky130_fd_sc_hd__decap_3 PHY_7227 ();
 sky130_fd_sc_hd__decap_3 PHY_7228 ();
 sky130_fd_sc_hd__decap_3 PHY_7229 ();
 sky130_fd_sc_hd__decap_3 PHY_7230 ();
 sky130_fd_sc_hd__decap_3 PHY_7231 ();
 sky130_fd_sc_hd__decap_3 PHY_7232 ();
 sky130_fd_sc_hd__decap_3 PHY_7233 ();
 sky130_fd_sc_hd__decap_3 PHY_7234 ();
 sky130_fd_sc_hd__decap_3 PHY_7235 ();
 sky130_fd_sc_hd__decap_3 PHY_7236 ();
 sky130_fd_sc_hd__decap_3 PHY_7237 ();
 sky130_fd_sc_hd__decap_3 PHY_7238 ();
 sky130_fd_sc_hd__decap_3 PHY_7239 ();
 sky130_fd_sc_hd__decap_3 PHY_7240 ();
 sky130_fd_sc_hd__decap_3 PHY_7241 ();
 sky130_fd_sc_hd__decap_3 PHY_7242 ();
 sky130_fd_sc_hd__decap_3 PHY_7243 ();
 sky130_fd_sc_hd__decap_3 PHY_7244 ();
 sky130_fd_sc_hd__decap_3 PHY_7245 ();
 sky130_fd_sc_hd__decap_3 PHY_7246 ();
 sky130_fd_sc_hd__decap_3 PHY_7247 ();
 sky130_fd_sc_hd__decap_3 PHY_7248 ();
 sky130_fd_sc_hd__decap_3 PHY_7249 ();
 sky130_fd_sc_hd__decap_3 PHY_7250 ();
 sky130_fd_sc_hd__decap_3 PHY_7251 ();
 sky130_fd_sc_hd__decap_3 PHY_7252 ();
 sky130_fd_sc_hd__decap_3 PHY_7253 ();
 sky130_fd_sc_hd__decap_3 PHY_7254 ();
 sky130_fd_sc_hd__decap_3 PHY_7255 ();
 sky130_fd_sc_hd__decap_3 PHY_7256 ();
 sky130_fd_sc_hd__decap_3 PHY_7257 ();
 sky130_fd_sc_hd__decap_3 PHY_7258 ();
 sky130_fd_sc_hd__decap_3 PHY_7259 ();
 sky130_fd_sc_hd__decap_3 PHY_7260 ();
 sky130_fd_sc_hd__decap_3 PHY_7261 ();
 sky130_fd_sc_hd__decap_3 PHY_7262 ();
 sky130_fd_sc_hd__decap_3 PHY_7263 ();
 sky130_fd_sc_hd__decap_3 PHY_7264 ();
 sky130_fd_sc_hd__decap_3 PHY_7265 ();
 sky130_fd_sc_hd__decap_3 PHY_7266 ();
 sky130_fd_sc_hd__decap_3 PHY_7267 ();
 sky130_fd_sc_hd__decap_3 PHY_7268 ();
 sky130_fd_sc_hd__decap_3 PHY_7269 ();
 sky130_fd_sc_hd__decap_3 PHY_7270 ();
 sky130_fd_sc_hd__decap_3 PHY_7271 ();
 sky130_fd_sc_hd__decap_3 PHY_7272 ();
 sky130_fd_sc_hd__decap_3 PHY_7273 ();
 sky130_fd_sc_hd__decap_3 PHY_7274 ();
 sky130_fd_sc_hd__decap_3 PHY_7275 ();
 sky130_fd_sc_hd__decap_3 PHY_7276 ();
 sky130_fd_sc_hd__decap_3 PHY_7277 ();
 sky130_fd_sc_hd__decap_3 PHY_7278 ();
 sky130_fd_sc_hd__decap_3 PHY_7279 ();
 sky130_fd_sc_hd__decap_3 PHY_7280 ();
 sky130_fd_sc_hd__decap_3 PHY_7281 ();
 sky130_fd_sc_hd__decap_3 PHY_7282 ();
 sky130_fd_sc_hd__decap_3 PHY_7283 ();
 sky130_fd_sc_hd__decap_3 PHY_7284 ();
 sky130_fd_sc_hd__decap_3 PHY_7285 ();
 sky130_fd_sc_hd__decap_3 PHY_7286 ();
 sky130_fd_sc_hd__decap_3 PHY_7287 ();
 sky130_fd_sc_hd__decap_3 PHY_7288 ();
 sky130_fd_sc_hd__decap_3 PHY_7289 ();
 sky130_fd_sc_hd__decap_3 PHY_7290 ();
 sky130_fd_sc_hd__decap_3 PHY_7291 ();
 sky130_fd_sc_hd__decap_3 PHY_7292 ();
 sky130_fd_sc_hd__decap_3 PHY_7293 ();
 sky130_fd_sc_hd__decap_3 PHY_7294 ();
 sky130_fd_sc_hd__decap_3 PHY_7295 ();
 sky130_fd_sc_hd__decap_3 PHY_7296 ();
 sky130_fd_sc_hd__decap_3 PHY_7297 ();
 sky130_fd_sc_hd__decap_3 PHY_7298 ();
 sky130_fd_sc_hd__decap_3 PHY_7299 ();
 sky130_fd_sc_hd__decap_3 PHY_7300 ();
 sky130_fd_sc_hd__decap_3 PHY_7301 ();
 sky130_fd_sc_hd__decap_3 PHY_7302 ();
 sky130_fd_sc_hd__decap_3 PHY_7303 ();
 sky130_fd_sc_hd__decap_3 PHY_7304 ();
 sky130_fd_sc_hd__decap_3 PHY_7305 ();
 sky130_fd_sc_hd__decap_3 PHY_7306 ();
 sky130_fd_sc_hd__decap_3 PHY_7307 ();
 sky130_fd_sc_hd__decap_3 PHY_7308 ();
 sky130_fd_sc_hd__decap_3 PHY_7309 ();
 sky130_fd_sc_hd__decap_3 PHY_7310 ();
 sky130_fd_sc_hd__decap_3 PHY_7311 ();
 sky130_fd_sc_hd__decap_3 PHY_7312 ();
 sky130_fd_sc_hd__decap_3 PHY_7313 ();
 sky130_fd_sc_hd__decap_3 PHY_7314 ();
 sky130_fd_sc_hd__decap_3 PHY_7315 ();
 sky130_fd_sc_hd__decap_3 PHY_7316 ();
 sky130_fd_sc_hd__decap_3 PHY_7317 ();
 sky130_fd_sc_hd__decap_3 PHY_7318 ();
 sky130_fd_sc_hd__decap_3 PHY_7319 ();
 sky130_fd_sc_hd__decap_3 PHY_7320 ();
 sky130_fd_sc_hd__decap_3 PHY_7321 ();
 sky130_fd_sc_hd__decap_3 PHY_7322 ();
 sky130_fd_sc_hd__decap_3 PHY_7323 ();
 sky130_fd_sc_hd__decap_3 PHY_7324 ();
 sky130_fd_sc_hd__decap_3 PHY_7325 ();
 sky130_fd_sc_hd__decap_3 PHY_7326 ();
 sky130_fd_sc_hd__decap_3 PHY_7327 ();
 sky130_fd_sc_hd__decap_3 PHY_7328 ();
 sky130_fd_sc_hd__decap_3 PHY_7329 ();
 sky130_fd_sc_hd__decap_3 PHY_7330 ();
 sky130_fd_sc_hd__decap_3 PHY_7331 ();
 sky130_fd_sc_hd__decap_3 PHY_7332 ();
 sky130_fd_sc_hd__decap_3 PHY_7333 ();
 sky130_fd_sc_hd__decap_3 PHY_7334 ();
 sky130_fd_sc_hd__decap_3 PHY_7335 ();
 sky130_fd_sc_hd__decap_3 PHY_7336 ();
 sky130_fd_sc_hd__decap_3 PHY_7337 ();
 sky130_fd_sc_hd__decap_3 PHY_7338 ();
 sky130_fd_sc_hd__decap_3 PHY_7339 ();
 sky130_fd_sc_hd__decap_3 PHY_7340 ();
 sky130_fd_sc_hd__decap_3 PHY_7341 ();
 sky130_fd_sc_hd__decap_3 PHY_7342 ();
 sky130_fd_sc_hd__decap_3 PHY_7343 ();
 sky130_fd_sc_hd__decap_3 PHY_7344 ();
 sky130_fd_sc_hd__decap_3 PHY_7345 ();
 sky130_fd_sc_hd__decap_3 PHY_7346 ();
 sky130_fd_sc_hd__decap_3 PHY_7347 ();
 sky130_fd_sc_hd__decap_3 PHY_7348 ();
 sky130_fd_sc_hd__decap_3 PHY_7349 ();
 sky130_fd_sc_hd__decap_3 PHY_7350 ();
 sky130_fd_sc_hd__decap_3 PHY_7351 ();
 sky130_fd_sc_hd__decap_3 PHY_7352 ();
 sky130_fd_sc_hd__decap_3 PHY_7353 ();
 sky130_fd_sc_hd__decap_3 PHY_7354 ();
 sky130_fd_sc_hd__decap_3 PHY_7355 ();
 sky130_fd_sc_hd__decap_3 PHY_7356 ();
 sky130_fd_sc_hd__decap_3 PHY_7357 ();
 sky130_fd_sc_hd__decap_3 PHY_7358 ();
 sky130_fd_sc_hd__decap_3 PHY_7359 ();
 sky130_fd_sc_hd__decap_3 PHY_7360 ();
 sky130_fd_sc_hd__decap_3 PHY_7361 ();
 sky130_fd_sc_hd__decap_3 PHY_7362 ();
 sky130_fd_sc_hd__decap_3 PHY_7363 ();
 sky130_fd_sc_hd__decap_3 PHY_7364 ();
 sky130_fd_sc_hd__decap_3 PHY_7365 ();
 sky130_fd_sc_hd__decap_3 PHY_7366 ();
 sky130_fd_sc_hd__decap_3 PHY_7367 ();
 sky130_fd_sc_hd__decap_3 PHY_7368 ();
 sky130_fd_sc_hd__decap_3 PHY_7369 ();
 sky130_fd_sc_hd__decap_3 PHY_7370 ();
 sky130_fd_sc_hd__decap_3 PHY_7371 ();
 sky130_fd_sc_hd__decap_3 PHY_7372 ();
 sky130_fd_sc_hd__decap_3 PHY_7373 ();
 sky130_fd_sc_hd__decap_3 PHY_7374 ();
 sky130_fd_sc_hd__decap_3 PHY_7375 ();
 sky130_fd_sc_hd__decap_3 PHY_7376 ();
 sky130_fd_sc_hd__decap_3 PHY_7377 ();
 sky130_fd_sc_hd__decap_3 PHY_7378 ();
 sky130_fd_sc_hd__decap_3 PHY_7379 ();
 sky130_fd_sc_hd__decap_3 PHY_7380 ();
 sky130_fd_sc_hd__decap_3 PHY_7381 ();
 sky130_fd_sc_hd__decap_3 PHY_7382 ();
 sky130_fd_sc_hd__decap_3 PHY_7383 ();
 sky130_fd_sc_hd__decap_3 PHY_7384 ();
 sky130_fd_sc_hd__decap_3 PHY_7385 ();
 sky130_fd_sc_hd__decap_3 PHY_7386 ();
 sky130_fd_sc_hd__decap_3 PHY_7387 ();
 sky130_fd_sc_hd__decap_3 PHY_7388 ();
 sky130_fd_sc_hd__decap_3 PHY_7389 ();
 sky130_fd_sc_hd__decap_3 PHY_7390 ();
 sky130_fd_sc_hd__decap_3 PHY_7391 ();
 sky130_fd_sc_hd__decap_3 PHY_7392 ();
 sky130_fd_sc_hd__decap_3 PHY_7393 ();
 sky130_fd_sc_hd__decap_3 PHY_7394 ();
 sky130_fd_sc_hd__decap_3 PHY_7395 ();
 sky130_fd_sc_hd__decap_3 PHY_7396 ();
 sky130_fd_sc_hd__decap_3 PHY_7397 ();
 sky130_fd_sc_hd__decap_3 PHY_7398 ();
 sky130_fd_sc_hd__decap_3 PHY_7399 ();
 sky130_fd_sc_hd__decap_3 PHY_7400 ();
 sky130_fd_sc_hd__decap_3 PHY_7401 ();
 sky130_fd_sc_hd__decap_3 PHY_7402 ();
 sky130_fd_sc_hd__decap_3 PHY_7403 ();
 sky130_fd_sc_hd__decap_3 PHY_7404 ();
 sky130_fd_sc_hd__decap_3 PHY_7405 ();
 sky130_fd_sc_hd__decap_3 PHY_7406 ();
 sky130_fd_sc_hd__decap_3 PHY_7407 ();
 sky130_fd_sc_hd__decap_3 PHY_7408 ();
 sky130_fd_sc_hd__decap_3 PHY_7409 ();
 sky130_fd_sc_hd__decap_3 PHY_7410 ();
 sky130_fd_sc_hd__decap_3 PHY_7411 ();
 sky130_fd_sc_hd__decap_3 PHY_7412 ();
 sky130_fd_sc_hd__decap_3 PHY_7413 ();
 sky130_fd_sc_hd__decap_3 PHY_7414 ();
 sky130_fd_sc_hd__decap_3 PHY_7415 ();
 sky130_fd_sc_hd__decap_3 PHY_7416 ();
 sky130_fd_sc_hd__decap_3 PHY_7417 ();
 sky130_fd_sc_hd__decap_3 PHY_7418 ();
 sky130_fd_sc_hd__decap_3 PHY_7419 ();
 sky130_fd_sc_hd__decap_3 PHY_7420 ();
 sky130_fd_sc_hd__decap_3 PHY_7421 ();
 sky130_fd_sc_hd__decap_3 PHY_7422 ();
 sky130_fd_sc_hd__decap_3 PHY_7423 ();
 sky130_fd_sc_hd__decap_3 PHY_7424 ();
 sky130_fd_sc_hd__decap_3 PHY_7425 ();
 sky130_fd_sc_hd__decap_3 PHY_7426 ();
 sky130_fd_sc_hd__decap_3 PHY_7427 ();
 sky130_fd_sc_hd__decap_3 PHY_7428 ();
 sky130_fd_sc_hd__decap_3 PHY_7429 ();
 sky130_fd_sc_hd__decap_3 PHY_7430 ();
 sky130_fd_sc_hd__decap_3 PHY_7431 ();
 sky130_fd_sc_hd__decap_3 PHY_7432 ();
 sky130_fd_sc_hd__decap_3 PHY_7433 ();
 sky130_fd_sc_hd__decap_3 PHY_7434 ();
 sky130_fd_sc_hd__decap_3 PHY_7435 ();
 sky130_fd_sc_hd__decap_3 PHY_7436 ();
 sky130_fd_sc_hd__decap_3 PHY_7437 ();
 sky130_fd_sc_hd__decap_3 PHY_7438 ();
 sky130_fd_sc_hd__decap_3 PHY_7439 ();
 sky130_fd_sc_hd__decap_3 PHY_7440 ();
 sky130_fd_sc_hd__decap_3 PHY_7441 ();
 sky130_fd_sc_hd__decap_3 PHY_7442 ();
 sky130_fd_sc_hd__decap_3 PHY_7443 ();
 sky130_fd_sc_hd__decap_3 PHY_7444 ();
 sky130_fd_sc_hd__decap_3 PHY_7445 ();
 sky130_fd_sc_hd__decap_3 PHY_7446 ();
 sky130_fd_sc_hd__decap_3 PHY_7447 ();
 sky130_fd_sc_hd__decap_3 PHY_7448 ();
 sky130_fd_sc_hd__decap_3 PHY_7449 ();
 sky130_fd_sc_hd__decap_3 PHY_7450 ();
 sky130_fd_sc_hd__decap_3 PHY_7451 ();
 sky130_fd_sc_hd__decap_3 PHY_7452 ();
 sky130_fd_sc_hd__decap_3 PHY_7453 ();
 sky130_fd_sc_hd__decap_3 PHY_7454 ();
 sky130_fd_sc_hd__decap_3 PHY_7455 ();
 sky130_fd_sc_hd__decap_3 PHY_7456 ();
 sky130_fd_sc_hd__decap_3 PHY_7457 ();
 sky130_fd_sc_hd__decap_3 PHY_7458 ();
 sky130_fd_sc_hd__decap_3 PHY_7459 ();
 sky130_fd_sc_hd__decap_3 PHY_7460 ();
 sky130_fd_sc_hd__decap_3 PHY_7461 ();
 sky130_fd_sc_hd__decap_3 PHY_7462 ();
 sky130_fd_sc_hd__decap_3 PHY_7463 ();
 sky130_fd_sc_hd__decap_3 PHY_7464 ();
 sky130_fd_sc_hd__decap_3 PHY_7465 ();
 sky130_fd_sc_hd__decap_3 PHY_7466 ();
 sky130_fd_sc_hd__decap_3 PHY_7467 ();
 sky130_fd_sc_hd__decap_3 PHY_7468 ();
 sky130_fd_sc_hd__decap_3 PHY_7469 ();
 sky130_fd_sc_hd__decap_3 PHY_7470 ();
 sky130_fd_sc_hd__decap_3 PHY_7471 ();
 sky130_fd_sc_hd__decap_3 PHY_7472 ();
 sky130_fd_sc_hd__decap_3 PHY_7473 ();
 sky130_fd_sc_hd__decap_3 PHY_7474 ();
 sky130_fd_sc_hd__decap_3 PHY_7475 ();
 sky130_fd_sc_hd__decap_3 PHY_7476 ();
 sky130_fd_sc_hd__decap_3 PHY_7477 ();
 sky130_fd_sc_hd__decap_3 PHY_7478 ();
 sky130_fd_sc_hd__decap_3 PHY_7479 ();
 sky130_fd_sc_hd__decap_3 PHY_7480 ();
 sky130_fd_sc_hd__decap_3 PHY_7481 ();
 sky130_fd_sc_hd__decap_3 PHY_7482 ();
 sky130_fd_sc_hd__decap_3 PHY_7483 ();
 sky130_fd_sc_hd__decap_3 PHY_7484 ();
 sky130_fd_sc_hd__decap_3 PHY_7485 ();
 sky130_fd_sc_hd__decap_3 PHY_7486 ();
 sky130_fd_sc_hd__decap_3 PHY_7487 ();
 sky130_fd_sc_hd__decap_3 PHY_7488 ();
 sky130_fd_sc_hd__decap_3 PHY_7489 ();
 sky130_fd_sc_hd__decap_3 PHY_7490 ();
 sky130_fd_sc_hd__decap_3 PHY_7491 ();
 sky130_fd_sc_hd__decap_3 PHY_7492 ();
 sky130_fd_sc_hd__decap_3 PHY_7493 ();
 sky130_fd_sc_hd__decap_3 PHY_7494 ();
 sky130_fd_sc_hd__decap_3 PHY_7495 ();
 sky130_fd_sc_hd__decap_3 PHY_7496 ();
 sky130_fd_sc_hd__decap_3 PHY_7497 ();
 sky130_fd_sc_hd__decap_3 PHY_7498 ();
 sky130_fd_sc_hd__decap_3 PHY_7499 ();
 sky130_fd_sc_hd__decap_3 PHY_7500 ();
 sky130_fd_sc_hd__decap_3 PHY_7501 ();
 sky130_fd_sc_hd__decap_3 PHY_7502 ();
 sky130_fd_sc_hd__decap_3 PHY_7503 ();
 sky130_fd_sc_hd__decap_3 PHY_7504 ();
 sky130_fd_sc_hd__decap_3 PHY_7505 ();
 sky130_fd_sc_hd__decap_3 PHY_7506 ();
 sky130_fd_sc_hd__decap_3 PHY_7507 ();
 sky130_fd_sc_hd__decap_3 PHY_7508 ();
 sky130_fd_sc_hd__decap_3 PHY_7509 ();
 sky130_fd_sc_hd__decap_3 PHY_7510 ();
 sky130_fd_sc_hd__decap_3 PHY_7511 ();
 sky130_fd_sc_hd__decap_3 PHY_7512 ();
 sky130_fd_sc_hd__decap_3 PHY_7513 ();
 sky130_fd_sc_hd__decap_3 PHY_7514 ();
 sky130_fd_sc_hd__decap_3 PHY_7515 ();
 sky130_fd_sc_hd__decap_3 PHY_7516 ();
 sky130_fd_sc_hd__decap_3 PHY_7517 ();
 sky130_fd_sc_hd__decap_3 PHY_7518 ();
 sky130_fd_sc_hd__decap_3 PHY_7519 ();
 sky130_fd_sc_hd__decap_3 PHY_7520 ();
 sky130_fd_sc_hd__decap_3 PHY_7521 ();
 sky130_fd_sc_hd__decap_3 PHY_7522 ();
 sky130_fd_sc_hd__decap_3 PHY_7523 ();
 sky130_fd_sc_hd__decap_3 PHY_7524 ();
 sky130_fd_sc_hd__decap_3 PHY_7525 ();
 sky130_fd_sc_hd__decap_3 PHY_7526 ();
 sky130_fd_sc_hd__decap_3 PHY_7527 ();
 sky130_fd_sc_hd__decap_3 PHY_7528 ();
 sky130_fd_sc_hd__decap_3 PHY_7529 ();
 sky130_fd_sc_hd__decap_3 PHY_7530 ();
 sky130_fd_sc_hd__decap_3 PHY_7531 ();
 sky130_fd_sc_hd__decap_3 PHY_7532 ();
 sky130_fd_sc_hd__decap_3 PHY_7533 ();
 sky130_fd_sc_hd__decap_3 PHY_7534 ();
 sky130_fd_sc_hd__decap_3 PHY_7535 ();
 sky130_fd_sc_hd__decap_3 PHY_7536 ();
 sky130_fd_sc_hd__decap_3 PHY_7537 ();
 sky130_fd_sc_hd__decap_3 PHY_7538 ();
 sky130_fd_sc_hd__decap_3 PHY_7539 ();
 sky130_fd_sc_hd__decap_3 PHY_7540 ();
 sky130_fd_sc_hd__decap_3 PHY_7541 ();
 sky130_fd_sc_hd__decap_3 PHY_7542 ();
 sky130_fd_sc_hd__decap_3 PHY_7543 ();
 sky130_fd_sc_hd__decap_3 PHY_7544 ();
 sky130_fd_sc_hd__decap_3 PHY_7545 ();
 sky130_fd_sc_hd__decap_3 PHY_7546 ();
 sky130_fd_sc_hd__decap_3 PHY_7547 ();
 sky130_fd_sc_hd__decap_3 PHY_7548 ();
 sky130_fd_sc_hd__decap_3 PHY_7549 ();
 sky130_fd_sc_hd__decap_3 PHY_7550 ();
 sky130_fd_sc_hd__decap_3 PHY_7551 ();
 sky130_fd_sc_hd__decap_3 PHY_7552 ();
 sky130_fd_sc_hd__decap_3 PHY_7553 ();
 sky130_fd_sc_hd__decap_3 PHY_7554 ();
 sky130_fd_sc_hd__decap_3 PHY_7555 ();
 sky130_fd_sc_hd__decap_3 PHY_7556 ();
 sky130_fd_sc_hd__decap_3 PHY_7557 ();
 sky130_fd_sc_hd__decap_3 PHY_7558 ();
 sky130_fd_sc_hd__decap_3 PHY_7559 ();
 sky130_fd_sc_hd__decap_3 PHY_7560 ();
 sky130_fd_sc_hd__decap_3 PHY_7561 ();
 sky130_fd_sc_hd__decap_3 PHY_7562 ();
 sky130_fd_sc_hd__decap_3 PHY_7563 ();
 sky130_fd_sc_hd__decap_3 PHY_7564 ();
 sky130_fd_sc_hd__decap_3 PHY_7565 ();
 sky130_fd_sc_hd__decap_3 PHY_7566 ();
 sky130_fd_sc_hd__decap_3 PHY_7567 ();
 sky130_fd_sc_hd__decap_3 PHY_7568 ();
 sky130_fd_sc_hd__decap_3 PHY_7569 ();
 sky130_fd_sc_hd__decap_3 PHY_7570 ();
 sky130_fd_sc_hd__decap_3 PHY_7571 ();
 sky130_fd_sc_hd__decap_3 PHY_7572 ();
 sky130_fd_sc_hd__decap_3 PHY_7573 ();
 sky130_fd_sc_hd__decap_3 PHY_7574 ();
 sky130_fd_sc_hd__decap_3 PHY_7575 ();
 sky130_fd_sc_hd__decap_3 PHY_7576 ();
 sky130_fd_sc_hd__decap_3 PHY_7577 ();
 sky130_fd_sc_hd__decap_3 PHY_7578 ();
 sky130_fd_sc_hd__decap_3 PHY_7579 ();
 sky130_fd_sc_hd__decap_3 PHY_7580 ();
 sky130_fd_sc_hd__decap_3 PHY_7581 ();
 sky130_fd_sc_hd__decap_3 PHY_7582 ();
 sky130_fd_sc_hd__decap_3 PHY_7583 ();
 sky130_fd_sc_hd__decap_3 PHY_7584 ();
 sky130_fd_sc_hd__decap_3 PHY_7585 ();
 sky130_fd_sc_hd__decap_3 PHY_7586 ();
 sky130_fd_sc_hd__decap_3 PHY_7587 ();
 sky130_fd_sc_hd__decap_3 PHY_7588 ();
 sky130_fd_sc_hd__decap_3 PHY_7589 ();
 sky130_fd_sc_hd__decap_3 PHY_7590 ();
 sky130_fd_sc_hd__decap_3 PHY_7591 ();
 sky130_fd_sc_hd__decap_3 PHY_7592 ();
 sky130_fd_sc_hd__decap_3 PHY_7593 ();
 sky130_fd_sc_hd__decap_3 PHY_7594 ();
 sky130_fd_sc_hd__decap_3 PHY_7595 ();
 sky130_fd_sc_hd__decap_3 PHY_7596 ();
 sky130_fd_sc_hd__decap_3 PHY_7597 ();
 sky130_fd_sc_hd__decap_3 PHY_7598 ();
 sky130_fd_sc_hd__decap_3 PHY_7599 ();
 sky130_fd_sc_hd__decap_3 PHY_7600 ();
 sky130_fd_sc_hd__decap_3 PHY_7601 ();
 sky130_fd_sc_hd__decap_3 PHY_7602 ();
 sky130_fd_sc_hd__decap_3 PHY_7603 ();
 sky130_fd_sc_hd__decap_3 PHY_7604 ();
 sky130_fd_sc_hd__decap_3 PHY_7605 ();
 sky130_fd_sc_hd__decap_3 PHY_7606 ();
 sky130_fd_sc_hd__decap_3 PHY_7607 ();
 sky130_fd_sc_hd__decap_3 PHY_7608 ();
 sky130_fd_sc_hd__decap_3 PHY_7609 ();
 sky130_fd_sc_hd__decap_3 PHY_7610 ();
 sky130_fd_sc_hd__decap_3 PHY_7611 ();
 sky130_fd_sc_hd__decap_3 PHY_7612 ();
 sky130_fd_sc_hd__decap_3 PHY_7613 ();
 sky130_fd_sc_hd__decap_3 PHY_7614 ();
 sky130_fd_sc_hd__decap_3 PHY_7615 ();
 sky130_fd_sc_hd__decap_3 PHY_7616 ();
 sky130_fd_sc_hd__decap_3 PHY_7617 ();
 sky130_fd_sc_hd__decap_3 PHY_7618 ();
 sky130_fd_sc_hd__decap_3 PHY_7619 ();
 sky130_fd_sc_hd__decap_3 PHY_7620 ();
 sky130_fd_sc_hd__decap_3 PHY_7621 ();
 sky130_fd_sc_hd__decap_3 PHY_7622 ();
 sky130_fd_sc_hd__decap_3 PHY_7623 ();
 sky130_fd_sc_hd__decap_3 PHY_7624 ();
 sky130_fd_sc_hd__decap_3 PHY_7625 ();
 sky130_fd_sc_hd__decap_3 PHY_7626 ();
 sky130_fd_sc_hd__decap_3 PHY_7627 ();
 sky130_fd_sc_hd__decap_3 PHY_7628 ();
 sky130_fd_sc_hd__decap_3 PHY_7629 ();
 sky130_fd_sc_hd__decap_3 PHY_7630 ();
 sky130_fd_sc_hd__decap_3 PHY_7631 ();
 sky130_fd_sc_hd__decap_3 PHY_7632 ();
 sky130_fd_sc_hd__decap_3 PHY_7633 ();
 sky130_fd_sc_hd__decap_3 PHY_7634 ();
 sky130_fd_sc_hd__decap_3 PHY_7635 ();
 sky130_fd_sc_hd__decap_3 PHY_7636 ();
 sky130_fd_sc_hd__decap_3 PHY_7637 ();
 sky130_fd_sc_hd__decap_3 PHY_7638 ();
 sky130_fd_sc_hd__decap_3 PHY_7639 ();
 sky130_fd_sc_hd__decap_3 PHY_7640 ();
 sky130_fd_sc_hd__decap_3 PHY_7641 ();
 sky130_fd_sc_hd__decap_3 PHY_7642 ();
 sky130_fd_sc_hd__decap_3 PHY_7643 ();
 sky130_fd_sc_hd__decap_3 PHY_7644 ();
 sky130_fd_sc_hd__decap_3 PHY_7645 ();
 sky130_fd_sc_hd__decap_3 PHY_7646 ();
 sky130_fd_sc_hd__decap_3 PHY_7647 ();
 sky130_fd_sc_hd__decap_3 PHY_7648 ();
 sky130_fd_sc_hd__decap_3 PHY_7649 ();
 sky130_fd_sc_hd__decap_3 PHY_7650 ();
 sky130_fd_sc_hd__decap_3 PHY_7651 ();
 sky130_fd_sc_hd__decap_3 PHY_7652 ();
 sky130_fd_sc_hd__decap_3 PHY_7653 ();
 sky130_fd_sc_hd__decap_3 PHY_7654 ();
 sky130_fd_sc_hd__decap_3 PHY_7655 ();
 sky130_fd_sc_hd__decap_3 PHY_7656 ();
 sky130_fd_sc_hd__decap_3 PHY_7657 ();
 sky130_fd_sc_hd__decap_3 PHY_7658 ();
 sky130_fd_sc_hd__decap_3 PHY_7659 ();
 sky130_fd_sc_hd__decap_3 PHY_7660 ();
 sky130_fd_sc_hd__decap_3 PHY_7661 ();
 sky130_fd_sc_hd__decap_3 PHY_7662 ();
 sky130_fd_sc_hd__decap_3 PHY_7663 ();
 sky130_fd_sc_hd__decap_3 PHY_7664 ();
 sky130_fd_sc_hd__decap_3 PHY_7665 ();
 sky130_fd_sc_hd__decap_3 PHY_7666 ();
 sky130_fd_sc_hd__decap_3 PHY_7667 ();
 sky130_fd_sc_hd__decap_3 PHY_7668 ();
 sky130_fd_sc_hd__decap_3 PHY_7669 ();
 sky130_fd_sc_hd__decap_3 PHY_7670 ();
 sky130_fd_sc_hd__decap_3 PHY_7671 ();
 sky130_fd_sc_hd__decap_3 PHY_7672 ();
 sky130_fd_sc_hd__decap_3 PHY_7673 ();
 sky130_fd_sc_hd__decap_3 PHY_7674 ();
 sky130_fd_sc_hd__decap_3 PHY_7675 ();
 sky130_fd_sc_hd__decap_3 PHY_7676 ();
 sky130_fd_sc_hd__decap_3 PHY_7677 ();
 sky130_fd_sc_hd__decap_3 PHY_7678 ();
 sky130_fd_sc_hd__decap_3 PHY_7679 ();
 sky130_fd_sc_hd__decap_3 PHY_7680 ();
 sky130_fd_sc_hd__decap_3 PHY_7681 ();
 sky130_fd_sc_hd__decap_3 PHY_7682 ();
 sky130_fd_sc_hd__decap_3 PHY_7683 ();
 sky130_fd_sc_hd__decap_3 PHY_7684 ();
 sky130_fd_sc_hd__decap_3 PHY_7685 ();
 sky130_fd_sc_hd__decap_3 PHY_7686 ();
 sky130_fd_sc_hd__decap_3 PHY_7687 ();
 sky130_fd_sc_hd__decap_3 PHY_7688 ();
 sky130_fd_sc_hd__decap_3 PHY_7689 ();
 sky130_fd_sc_hd__decap_3 PHY_7690 ();
 sky130_fd_sc_hd__decap_3 PHY_7691 ();
 sky130_fd_sc_hd__decap_3 PHY_7692 ();
 sky130_fd_sc_hd__decap_3 PHY_7693 ();
 sky130_fd_sc_hd__decap_3 PHY_7694 ();
 sky130_fd_sc_hd__decap_3 PHY_7695 ();
 sky130_fd_sc_hd__decap_3 PHY_7696 ();
 sky130_fd_sc_hd__decap_3 PHY_7697 ();
 sky130_fd_sc_hd__decap_3 PHY_7698 ();
 sky130_fd_sc_hd__decap_3 PHY_7699 ();
 sky130_fd_sc_hd__decap_3 PHY_7700 ();
 sky130_fd_sc_hd__decap_3 PHY_7701 ();
 sky130_fd_sc_hd__decap_3 PHY_7702 ();
 sky130_fd_sc_hd__decap_3 PHY_7703 ();
 sky130_fd_sc_hd__decap_3 PHY_7704 ();
 sky130_fd_sc_hd__decap_3 PHY_7705 ();
 sky130_fd_sc_hd__decap_3 PHY_7706 ();
 sky130_fd_sc_hd__decap_3 PHY_7707 ();
 sky130_fd_sc_hd__decap_3 PHY_7708 ();
 sky130_fd_sc_hd__decap_3 PHY_7709 ();
 sky130_fd_sc_hd__decap_3 PHY_7710 ();
 sky130_fd_sc_hd__decap_3 PHY_7711 ();
 sky130_fd_sc_hd__decap_3 PHY_7712 ();
 sky130_fd_sc_hd__decap_3 PHY_7713 ();
 sky130_fd_sc_hd__decap_3 PHY_7714 ();
 sky130_fd_sc_hd__decap_3 PHY_7715 ();
 sky130_fd_sc_hd__decap_3 PHY_7716 ();
 sky130_fd_sc_hd__decap_3 PHY_7717 ();
 sky130_fd_sc_hd__decap_3 PHY_7718 ();
 sky130_fd_sc_hd__decap_3 PHY_7719 ();
 sky130_fd_sc_hd__decap_3 PHY_7720 ();
 sky130_fd_sc_hd__decap_3 PHY_7721 ();
 sky130_fd_sc_hd__decap_3 PHY_7722 ();
 sky130_fd_sc_hd__decap_3 PHY_7723 ();
 sky130_fd_sc_hd__decap_3 PHY_7724 ();
 sky130_fd_sc_hd__decap_3 PHY_7725 ();
 sky130_fd_sc_hd__decap_3 PHY_7726 ();
 sky130_fd_sc_hd__decap_3 PHY_7727 ();
 sky130_fd_sc_hd__decap_3 PHY_7728 ();
 sky130_fd_sc_hd__decap_3 PHY_7729 ();
 sky130_fd_sc_hd__decap_3 PHY_7730 ();
 sky130_fd_sc_hd__decap_3 PHY_7731 ();
 sky130_fd_sc_hd__decap_3 PHY_7732 ();
 sky130_fd_sc_hd__decap_3 PHY_7733 ();
 sky130_fd_sc_hd__decap_3 PHY_7734 ();
 sky130_fd_sc_hd__decap_3 PHY_7735 ();
 sky130_fd_sc_hd__decap_3 PHY_7736 ();
 sky130_fd_sc_hd__decap_3 PHY_7737 ();
 sky130_fd_sc_hd__decap_3 PHY_7738 ();
 sky130_fd_sc_hd__decap_3 PHY_7739 ();
 sky130_fd_sc_hd__decap_3 PHY_7740 ();
 sky130_fd_sc_hd__decap_3 PHY_7741 ();
 sky130_fd_sc_hd__decap_3 PHY_7742 ();
 sky130_fd_sc_hd__decap_3 PHY_7743 ();
 sky130_fd_sc_hd__decap_3 PHY_7744 ();
 sky130_fd_sc_hd__decap_3 PHY_7745 ();
 sky130_fd_sc_hd__decap_3 PHY_7746 ();
 sky130_fd_sc_hd__decap_3 PHY_7747 ();
 sky130_fd_sc_hd__decap_3 PHY_7748 ();
 sky130_fd_sc_hd__decap_3 PHY_7749 ();
 sky130_fd_sc_hd__decap_3 PHY_7750 ();
 sky130_fd_sc_hd__decap_3 PHY_7751 ();
 sky130_fd_sc_hd__decap_3 PHY_7752 ();
 sky130_fd_sc_hd__decap_3 PHY_7753 ();
 sky130_fd_sc_hd__decap_3 PHY_7754 ();
 sky130_fd_sc_hd__decap_3 PHY_7755 ();
 sky130_fd_sc_hd__decap_3 PHY_7756 ();
 sky130_fd_sc_hd__decap_3 PHY_7757 ();
 sky130_fd_sc_hd__decap_3 PHY_7758 ();
 sky130_fd_sc_hd__decap_3 PHY_7759 ();
 sky130_fd_sc_hd__decap_3 PHY_7760 ();
 sky130_fd_sc_hd__decap_3 PHY_7761 ();
 sky130_fd_sc_hd__decap_3 PHY_7762 ();
 sky130_fd_sc_hd__decap_3 PHY_7763 ();
 sky130_fd_sc_hd__decap_3 PHY_7764 ();
 sky130_fd_sc_hd__decap_3 PHY_7765 ();
 sky130_fd_sc_hd__decap_3 PHY_7766 ();
 sky130_fd_sc_hd__decap_3 PHY_7767 ();
 sky130_fd_sc_hd__decap_3 PHY_7768 ();
 sky130_fd_sc_hd__decap_3 PHY_7769 ();
 sky130_fd_sc_hd__decap_3 PHY_7770 ();
 sky130_fd_sc_hd__decap_3 PHY_7771 ();
 sky130_fd_sc_hd__decap_3 PHY_7772 ();
 sky130_fd_sc_hd__decap_3 PHY_7773 ();
 sky130_fd_sc_hd__decap_3 PHY_7774 ();
 sky130_fd_sc_hd__decap_3 PHY_7775 ();
 sky130_fd_sc_hd__decap_3 PHY_7776 ();
 sky130_fd_sc_hd__decap_3 PHY_7777 ();
 sky130_fd_sc_hd__decap_3 PHY_7778 ();
 sky130_fd_sc_hd__decap_3 PHY_7779 ();
 sky130_fd_sc_hd__decap_3 PHY_7780 ();
 sky130_fd_sc_hd__decap_3 PHY_7781 ();
 sky130_fd_sc_hd__decap_3 PHY_7782 ();
 sky130_fd_sc_hd__decap_3 PHY_7783 ();
 sky130_fd_sc_hd__decap_3 PHY_7784 ();
 sky130_fd_sc_hd__decap_3 PHY_7785 ();
 sky130_fd_sc_hd__decap_3 PHY_7786 ();
 sky130_fd_sc_hd__decap_3 PHY_7787 ();
 sky130_fd_sc_hd__decap_3 PHY_7788 ();
 sky130_fd_sc_hd__decap_3 PHY_7789 ();
 sky130_fd_sc_hd__decap_3 PHY_7790 ();
 sky130_fd_sc_hd__decap_3 PHY_7791 ();
 sky130_fd_sc_hd__decap_3 PHY_7792 ();
 sky130_fd_sc_hd__decap_3 PHY_7793 ();
 sky130_fd_sc_hd__decap_3 PHY_7794 ();
 sky130_fd_sc_hd__decap_3 PHY_7795 ();
 sky130_fd_sc_hd__decap_3 PHY_7796 ();
 sky130_fd_sc_hd__decap_3 PHY_7797 ();
 sky130_fd_sc_hd__decap_3 PHY_7798 ();
 sky130_fd_sc_hd__decap_3 PHY_7799 ();
 sky130_fd_sc_hd__decap_3 PHY_7800 ();
 sky130_fd_sc_hd__decap_3 PHY_7801 ();
 sky130_fd_sc_hd__decap_3 PHY_7802 ();
 sky130_fd_sc_hd__decap_3 PHY_7803 ();
 sky130_fd_sc_hd__decap_3 PHY_7804 ();
 sky130_fd_sc_hd__decap_3 PHY_7805 ();
 sky130_fd_sc_hd__decap_3 PHY_7806 ();
 sky130_fd_sc_hd__decap_3 PHY_7807 ();
 sky130_fd_sc_hd__decap_3 PHY_7808 ();
 sky130_fd_sc_hd__decap_3 PHY_7809 ();
 sky130_fd_sc_hd__decap_3 PHY_7810 ();
 sky130_fd_sc_hd__decap_3 PHY_7811 ();
 sky130_fd_sc_hd__decap_3 PHY_7812 ();
 sky130_fd_sc_hd__decap_3 PHY_7813 ();
 sky130_fd_sc_hd__decap_3 PHY_7814 ();
 sky130_fd_sc_hd__decap_3 PHY_7815 ();
 sky130_fd_sc_hd__decap_3 PHY_7816 ();
 sky130_fd_sc_hd__decap_3 PHY_7817 ();
 sky130_fd_sc_hd__decap_3 PHY_7818 ();
 sky130_fd_sc_hd__decap_3 PHY_7819 ();
 sky130_fd_sc_hd__decap_3 PHY_7820 ();
 sky130_fd_sc_hd__decap_3 PHY_7821 ();
 sky130_fd_sc_hd__decap_3 PHY_7822 ();
 sky130_fd_sc_hd__decap_3 PHY_7823 ();
 sky130_fd_sc_hd__decap_3 PHY_7824 ();
 sky130_fd_sc_hd__decap_3 PHY_7825 ();
 sky130_fd_sc_hd__decap_3 PHY_7826 ();
 sky130_fd_sc_hd__decap_3 PHY_7827 ();
 sky130_fd_sc_hd__decap_3 PHY_7828 ();
 sky130_fd_sc_hd__decap_3 PHY_7829 ();
 sky130_fd_sc_hd__decap_3 PHY_7830 ();
 sky130_fd_sc_hd__decap_3 PHY_7831 ();
 sky130_fd_sc_hd__decap_3 PHY_7832 ();
 sky130_fd_sc_hd__decap_3 PHY_7833 ();
 sky130_fd_sc_hd__decap_3 PHY_7834 ();
 sky130_fd_sc_hd__decap_3 PHY_7835 ();
 sky130_fd_sc_hd__decap_3 PHY_7836 ();
 sky130_fd_sc_hd__decap_3 PHY_7837 ();
 sky130_fd_sc_hd__decap_3 PHY_7838 ();
 sky130_fd_sc_hd__decap_3 PHY_7839 ();
 sky130_fd_sc_hd__decap_3 PHY_7840 ();
 sky130_fd_sc_hd__decap_3 PHY_7841 ();
 sky130_fd_sc_hd__decap_3 PHY_7842 ();
 sky130_fd_sc_hd__decap_3 PHY_7843 ();
 sky130_fd_sc_hd__decap_3 PHY_7844 ();
 sky130_fd_sc_hd__decap_3 PHY_7845 ();
 sky130_fd_sc_hd__decap_3 PHY_7846 ();
 sky130_fd_sc_hd__decap_3 PHY_7847 ();
 sky130_fd_sc_hd__decap_3 PHY_7848 ();
 sky130_fd_sc_hd__decap_3 PHY_7849 ();
 sky130_fd_sc_hd__decap_3 PHY_7850 ();
 sky130_fd_sc_hd__decap_3 PHY_7851 ();
 sky130_fd_sc_hd__decap_3 PHY_7852 ();
 sky130_fd_sc_hd__decap_3 PHY_7853 ();
 sky130_fd_sc_hd__decap_3 PHY_7854 ();
 sky130_fd_sc_hd__decap_3 PHY_7855 ();
 sky130_fd_sc_hd__decap_3 PHY_7856 ();
 sky130_fd_sc_hd__decap_3 PHY_7857 ();
 sky130_fd_sc_hd__decap_3 PHY_7858 ();
 sky130_fd_sc_hd__decap_3 PHY_7859 ();
 sky130_fd_sc_hd__decap_3 PHY_7860 ();
 sky130_fd_sc_hd__decap_3 PHY_7861 ();
 sky130_fd_sc_hd__decap_3 PHY_7862 ();
 sky130_fd_sc_hd__decap_3 PHY_7863 ();
 sky130_fd_sc_hd__decap_3 PHY_7864 ();
 sky130_fd_sc_hd__decap_3 PHY_7865 ();
 sky130_fd_sc_hd__decap_3 PHY_7866 ();
 sky130_fd_sc_hd__decap_3 PHY_7867 ();
 sky130_fd_sc_hd__decap_3 PHY_7868 ();
 sky130_fd_sc_hd__decap_3 PHY_7869 ();
 sky130_fd_sc_hd__decap_3 PHY_7870 ();
 sky130_fd_sc_hd__decap_3 PHY_7871 ();
 sky130_fd_sc_hd__decap_3 PHY_7872 ();
 sky130_fd_sc_hd__decap_3 PHY_7873 ();
 sky130_fd_sc_hd__decap_3 PHY_7874 ();
 sky130_fd_sc_hd__decap_3 PHY_7875 ();
 sky130_fd_sc_hd__decap_3 PHY_7876 ();
 sky130_fd_sc_hd__decap_3 PHY_7877 ();
 sky130_fd_sc_hd__decap_3 PHY_7878 ();
 sky130_fd_sc_hd__decap_3 PHY_7879 ();
 sky130_fd_sc_hd__decap_3 PHY_7880 ();
 sky130_fd_sc_hd__decap_3 PHY_7881 ();
 sky130_fd_sc_hd__decap_3 PHY_7882 ();
 sky130_fd_sc_hd__decap_3 PHY_7883 ();
 sky130_fd_sc_hd__decap_3 PHY_7884 ();
 sky130_fd_sc_hd__decap_3 PHY_7885 ();
 sky130_fd_sc_hd__decap_3 PHY_7886 ();
 sky130_fd_sc_hd__decap_3 PHY_7887 ();
 sky130_fd_sc_hd__decap_3 PHY_7888 ();
 sky130_fd_sc_hd__decap_3 PHY_7889 ();
 sky130_fd_sc_hd__decap_3 PHY_7890 ();
 sky130_fd_sc_hd__decap_3 PHY_7891 ();
 sky130_fd_sc_hd__decap_3 PHY_7892 ();
 sky130_fd_sc_hd__decap_3 PHY_7893 ();
 sky130_fd_sc_hd__decap_3 PHY_7894 ();
 sky130_fd_sc_hd__decap_3 PHY_7895 ();
 sky130_fd_sc_hd__decap_3 PHY_7896 ();
 sky130_fd_sc_hd__decap_3 PHY_7897 ();
 sky130_fd_sc_hd__decap_3 PHY_7898 ();
 sky130_fd_sc_hd__decap_3 PHY_7899 ();
 sky130_fd_sc_hd__decap_3 PHY_7900 ();
 sky130_fd_sc_hd__decap_3 PHY_7901 ();
 sky130_fd_sc_hd__decap_3 PHY_7902 ();
 sky130_fd_sc_hd__decap_3 PHY_7903 ();
 sky130_fd_sc_hd__decap_3 PHY_7904 ();
 sky130_fd_sc_hd__decap_3 PHY_7905 ();
 sky130_fd_sc_hd__decap_3 PHY_7906 ();
 sky130_fd_sc_hd__decap_3 PHY_7907 ();
 sky130_fd_sc_hd__decap_3 PHY_7908 ();
 sky130_fd_sc_hd__decap_3 PHY_7909 ();
 sky130_fd_sc_hd__decap_3 PHY_7910 ();
 sky130_fd_sc_hd__decap_3 PHY_7911 ();
 sky130_fd_sc_hd__decap_3 PHY_7912 ();
 sky130_fd_sc_hd__decap_3 PHY_7913 ();
 sky130_fd_sc_hd__decap_3 PHY_7914 ();
 sky130_fd_sc_hd__decap_3 PHY_7915 ();
 sky130_fd_sc_hd__decap_3 PHY_7916 ();
 sky130_fd_sc_hd__decap_3 PHY_7917 ();
 sky130_fd_sc_hd__decap_3 PHY_7918 ();
 sky130_fd_sc_hd__decap_3 PHY_7919 ();
 sky130_fd_sc_hd__decap_3 PHY_7920 ();
 sky130_fd_sc_hd__decap_3 PHY_7921 ();
 sky130_fd_sc_hd__decap_3 PHY_7922 ();
 sky130_fd_sc_hd__decap_3 PHY_7923 ();
 sky130_fd_sc_hd__decap_3 PHY_7924 ();
 sky130_fd_sc_hd__decap_3 PHY_7925 ();
 sky130_fd_sc_hd__decap_3 PHY_7926 ();
 sky130_fd_sc_hd__decap_3 PHY_7927 ();
 sky130_fd_sc_hd__decap_3 PHY_7928 ();
 sky130_fd_sc_hd__decap_3 PHY_7929 ();
 sky130_fd_sc_hd__decap_3 PHY_7930 ();
 sky130_fd_sc_hd__decap_3 PHY_7931 ();
 sky130_fd_sc_hd__decap_3 PHY_7932 ();
 sky130_fd_sc_hd__decap_3 PHY_7933 ();
 sky130_fd_sc_hd__decap_3 PHY_7934 ();
 sky130_fd_sc_hd__decap_3 PHY_7935 ();
 sky130_fd_sc_hd__decap_3 PHY_7936 ();
 sky130_fd_sc_hd__decap_3 PHY_7937 ();
 sky130_fd_sc_hd__decap_3 PHY_7938 ();
 sky130_fd_sc_hd__decap_3 PHY_7939 ();
 sky130_fd_sc_hd__decap_3 PHY_7940 ();
 sky130_fd_sc_hd__decap_3 PHY_7941 ();
 sky130_fd_sc_hd__decap_3 PHY_7942 ();
 sky130_fd_sc_hd__decap_3 PHY_7943 ();
 sky130_fd_sc_hd__decap_3 PHY_7944 ();
 sky130_fd_sc_hd__decap_3 PHY_7945 ();
 sky130_fd_sc_hd__decap_3 PHY_7946 ();
 sky130_fd_sc_hd__decap_3 PHY_7947 ();
 sky130_fd_sc_hd__decap_3 PHY_7948 ();
 sky130_fd_sc_hd__decap_3 PHY_7949 ();
 sky130_fd_sc_hd__decap_3 PHY_7950 ();
 sky130_fd_sc_hd__decap_3 PHY_7951 ();
 sky130_fd_sc_hd__decap_3 PHY_7952 ();
 sky130_fd_sc_hd__decap_3 PHY_7953 ();
 sky130_fd_sc_hd__decap_3 PHY_7954 ();
 sky130_fd_sc_hd__decap_3 PHY_7955 ();
 sky130_fd_sc_hd__decap_3 PHY_7956 ();
 sky130_fd_sc_hd__decap_3 PHY_7957 ();
 sky130_fd_sc_hd__decap_3 PHY_7958 ();
 sky130_fd_sc_hd__decap_3 PHY_7959 ();
 sky130_fd_sc_hd__decap_3 PHY_7960 ();
 sky130_fd_sc_hd__decap_3 PHY_7961 ();
 sky130_fd_sc_hd__decap_3 PHY_7962 ();
 sky130_fd_sc_hd__decap_3 PHY_7963 ();
 sky130_fd_sc_hd__decap_3 PHY_7964 ();
 sky130_fd_sc_hd__decap_3 PHY_7965 ();
 sky130_fd_sc_hd__decap_3 PHY_7966 ();
 sky130_fd_sc_hd__decap_3 PHY_7967 ();
 sky130_fd_sc_hd__decap_3 PHY_7968 ();
 sky130_fd_sc_hd__decap_3 PHY_7969 ();
 sky130_fd_sc_hd__decap_3 PHY_7970 ();
 sky130_fd_sc_hd__decap_3 PHY_7971 ();
 sky130_fd_sc_hd__decap_3 PHY_7972 ();
 sky130_fd_sc_hd__decap_3 PHY_7973 ();
 sky130_fd_sc_hd__decap_3 PHY_7974 ();
 sky130_fd_sc_hd__decap_3 PHY_7975 ();
 sky130_fd_sc_hd__decap_3 PHY_7976 ();
 sky130_fd_sc_hd__decap_3 PHY_7977 ();
 sky130_fd_sc_hd__decap_3 PHY_7978 ();
 sky130_fd_sc_hd__decap_3 PHY_7979 ();
 sky130_fd_sc_hd__decap_3 PHY_7980 ();
 sky130_fd_sc_hd__decap_3 PHY_7981 ();
 sky130_fd_sc_hd__decap_3 PHY_7982 ();
 sky130_fd_sc_hd__decap_3 PHY_7983 ();
 sky130_fd_sc_hd__decap_3 PHY_7984 ();
 sky130_fd_sc_hd__decap_3 PHY_7985 ();
 sky130_fd_sc_hd__decap_3 PHY_7986 ();
 sky130_fd_sc_hd__decap_3 PHY_7987 ();
 sky130_fd_sc_hd__decap_3 PHY_7988 ();
 sky130_fd_sc_hd__decap_3 PHY_7989 ();
 sky130_fd_sc_hd__decap_3 PHY_7990 ();
 sky130_fd_sc_hd__decap_3 PHY_7991 ();
 sky130_fd_sc_hd__decap_3 PHY_7992 ();
 sky130_fd_sc_hd__decap_3 PHY_7993 ();
 sky130_fd_sc_hd__decap_3 PHY_7994 ();
 sky130_fd_sc_hd__decap_3 PHY_7995 ();
 sky130_fd_sc_hd__decap_3 PHY_7996 ();
 sky130_fd_sc_hd__decap_3 PHY_7997 ();
 sky130_fd_sc_hd__decap_3 PHY_7998 ();
 sky130_fd_sc_hd__decap_3 PHY_7999 ();
 sky130_fd_sc_hd__decap_3 PHY_8000 ();
 sky130_fd_sc_hd__decap_3 PHY_8001 ();
 sky130_fd_sc_hd__decap_3 PHY_8002 ();
 sky130_fd_sc_hd__decap_3 PHY_8003 ();
 sky130_fd_sc_hd__decap_3 PHY_8004 ();
 sky130_fd_sc_hd__decap_3 PHY_8005 ();
 sky130_fd_sc_hd__decap_3 PHY_8006 ();
 sky130_fd_sc_hd__decap_3 PHY_8007 ();
 sky130_fd_sc_hd__decap_3 PHY_8008 ();
 sky130_fd_sc_hd__decap_3 PHY_8009 ();
 sky130_fd_sc_hd__decap_3 PHY_8010 ();
 sky130_fd_sc_hd__decap_3 PHY_8011 ();
 sky130_fd_sc_hd__decap_3 PHY_8012 ();
 sky130_fd_sc_hd__decap_3 PHY_8013 ();
 sky130_fd_sc_hd__decap_3 PHY_8014 ();
 sky130_fd_sc_hd__decap_3 PHY_8015 ();
 sky130_fd_sc_hd__decap_3 PHY_8016 ();
 sky130_fd_sc_hd__decap_3 PHY_8017 ();
 sky130_fd_sc_hd__decap_3 PHY_8018 ();
 sky130_fd_sc_hd__decap_3 PHY_8019 ();
 sky130_fd_sc_hd__decap_3 PHY_8020 ();
 sky130_fd_sc_hd__decap_3 PHY_8021 ();
 sky130_fd_sc_hd__decap_3 PHY_8022 ();
 sky130_fd_sc_hd__decap_3 PHY_8023 ();
 sky130_fd_sc_hd__decap_3 PHY_8024 ();
 sky130_fd_sc_hd__decap_3 PHY_8025 ();
 sky130_fd_sc_hd__decap_3 PHY_8026 ();
 sky130_fd_sc_hd__decap_3 PHY_8027 ();
 sky130_fd_sc_hd__decap_3 PHY_8028 ();
 sky130_fd_sc_hd__decap_3 PHY_8029 ();
 sky130_fd_sc_hd__decap_3 PHY_8030 ();
 sky130_fd_sc_hd__decap_3 PHY_8031 ();
 sky130_fd_sc_hd__decap_3 PHY_8032 ();
 sky130_fd_sc_hd__decap_3 PHY_8033 ();
 sky130_fd_sc_hd__decap_3 PHY_8034 ();
 sky130_fd_sc_hd__decap_3 PHY_8035 ();
 sky130_fd_sc_hd__decap_3 PHY_8036 ();
 sky130_fd_sc_hd__decap_3 PHY_8037 ();
 sky130_fd_sc_hd__decap_3 PHY_8038 ();
 sky130_fd_sc_hd__decap_3 PHY_8039 ();
 sky130_fd_sc_hd__decap_3 PHY_8040 ();
 sky130_fd_sc_hd__decap_3 PHY_8041 ();
 sky130_fd_sc_hd__decap_3 PHY_8042 ();
 sky130_fd_sc_hd__decap_3 PHY_8043 ();
 sky130_fd_sc_hd__decap_3 PHY_8044 ();
 sky130_fd_sc_hd__decap_3 PHY_8045 ();
 sky130_fd_sc_hd__decap_3 PHY_8046 ();
 sky130_fd_sc_hd__decap_3 PHY_8047 ();
 sky130_fd_sc_hd__decap_3 PHY_8048 ();
 sky130_fd_sc_hd__decap_3 PHY_8049 ();
 sky130_fd_sc_hd__decap_3 PHY_8050 ();
 sky130_fd_sc_hd__decap_3 PHY_8051 ();
 sky130_fd_sc_hd__decap_3 PHY_8052 ();
 sky130_fd_sc_hd__decap_3 PHY_8053 ();
 sky130_fd_sc_hd__decap_3 PHY_8054 ();
 sky130_fd_sc_hd__decap_3 PHY_8055 ();
 sky130_fd_sc_hd__decap_3 PHY_8056 ();
 sky130_fd_sc_hd__decap_3 PHY_8057 ();
 sky130_fd_sc_hd__decap_3 PHY_8058 ();
 sky130_fd_sc_hd__decap_3 PHY_8059 ();
 sky130_fd_sc_hd__decap_3 PHY_8060 ();
 sky130_fd_sc_hd__decap_3 PHY_8061 ();
 sky130_fd_sc_hd__decap_3 PHY_8062 ();
 sky130_fd_sc_hd__decap_3 PHY_8063 ();
 sky130_fd_sc_hd__decap_3 PHY_8064 ();
 sky130_fd_sc_hd__decap_3 PHY_8065 ();
 sky130_fd_sc_hd__decap_3 PHY_8066 ();
 sky130_fd_sc_hd__decap_3 PHY_8067 ();
 sky130_fd_sc_hd__decap_3 PHY_8068 ();
 sky130_fd_sc_hd__decap_3 PHY_8069 ();
 sky130_fd_sc_hd__decap_3 PHY_8070 ();
 sky130_fd_sc_hd__decap_3 PHY_8071 ();
 sky130_fd_sc_hd__decap_3 PHY_8072 ();
 sky130_fd_sc_hd__decap_3 PHY_8073 ();
 sky130_fd_sc_hd__decap_3 PHY_8074 ();
 sky130_fd_sc_hd__decap_3 PHY_8075 ();
 sky130_fd_sc_hd__decap_3 PHY_8076 ();
 sky130_fd_sc_hd__decap_3 PHY_8077 ();
 sky130_fd_sc_hd__decap_3 PHY_8078 ();
 sky130_fd_sc_hd__decap_3 PHY_8079 ();
 sky130_fd_sc_hd__decap_3 PHY_8080 ();
 sky130_fd_sc_hd__decap_3 PHY_8081 ();
 sky130_fd_sc_hd__decap_3 PHY_8082 ();
 sky130_fd_sc_hd__decap_3 PHY_8083 ();
 sky130_fd_sc_hd__decap_3 PHY_8084 ();
 sky130_fd_sc_hd__decap_3 PHY_8085 ();
 sky130_fd_sc_hd__decap_3 PHY_8086 ();
 sky130_fd_sc_hd__decap_3 PHY_8087 ();
 sky130_fd_sc_hd__decap_3 PHY_8088 ();
 sky130_fd_sc_hd__decap_3 PHY_8089 ();
 sky130_fd_sc_hd__decap_3 PHY_8090 ();
 sky130_fd_sc_hd__decap_3 PHY_8091 ();
 sky130_fd_sc_hd__decap_3 PHY_8092 ();
 sky130_fd_sc_hd__decap_3 PHY_8093 ();
 sky130_fd_sc_hd__decap_3 PHY_8094 ();
 sky130_fd_sc_hd__decap_3 PHY_8095 ();
 sky130_fd_sc_hd__decap_3 PHY_8096 ();
 sky130_fd_sc_hd__decap_3 PHY_8097 ();
 sky130_fd_sc_hd__decap_3 PHY_8098 ();
 sky130_fd_sc_hd__decap_3 PHY_8099 ();
 sky130_fd_sc_hd__decap_3 PHY_8100 ();
 sky130_fd_sc_hd__decap_3 PHY_8101 ();
 sky130_fd_sc_hd__decap_3 PHY_8102 ();
 sky130_fd_sc_hd__decap_3 PHY_8103 ();
 sky130_fd_sc_hd__decap_3 PHY_8104 ();
 sky130_fd_sc_hd__decap_3 PHY_8105 ();
 sky130_fd_sc_hd__decap_3 PHY_8106 ();
 sky130_fd_sc_hd__decap_3 PHY_8107 ();
 sky130_fd_sc_hd__decap_3 PHY_8108 ();
 sky130_fd_sc_hd__decap_3 PHY_8109 ();
 sky130_fd_sc_hd__decap_3 PHY_8110 ();
 sky130_fd_sc_hd__decap_3 PHY_8111 ();
 sky130_fd_sc_hd__decap_3 PHY_8112 ();
 sky130_fd_sc_hd__decap_3 PHY_8113 ();
 sky130_fd_sc_hd__decap_3 PHY_8114 ();
 sky130_fd_sc_hd__decap_3 PHY_8115 ();
 sky130_fd_sc_hd__decap_3 PHY_8116 ();
 sky130_fd_sc_hd__decap_3 PHY_8117 ();
 sky130_fd_sc_hd__decap_3 PHY_8118 ();
 sky130_fd_sc_hd__decap_3 PHY_8119 ();
 sky130_fd_sc_hd__decap_3 PHY_8120 ();
 sky130_fd_sc_hd__decap_3 PHY_8121 ();
 sky130_fd_sc_hd__decap_3 PHY_8122 ();
 sky130_fd_sc_hd__decap_3 PHY_8123 ();
 sky130_fd_sc_hd__decap_3 PHY_8124 ();
 sky130_fd_sc_hd__decap_3 PHY_8125 ();
 sky130_fd_sc_hd__decap_3 PHY_8126 ();
 sky130_fd_sc_hd__decap_3 PHY_8127 ();
 sky130_fd_sc_hd__decap_3 PHY_8128 ();
 sky130_fd_sc_hd__decap_3 PHY_8129 ();
 sky130_fd_sc_hd__decap_3 PHY_8130 ();
 sky130_fd_sc_hd__decap_3 PHY_8131 ();
 sky130_fd_sc_hd__decap_3 PHY_8132 ();
 sky130_fd_sc_hd__decap_3 PHY_8133 ();
 sky130_fd_sc_hd__decap_3 PHY_8134 ();
 sky130_fd_sc_hd__decap_3 PHY_8135 ();
 sky130_fd_sc_hd__decap_3 PHY_8136 ();
 sky130_fd_sc_hd__decap_3 PHY_8137 ();
 sky130_fd_sc_hd__decap_3 PHY_8138 ();
 sky130_fd_sc_hd__decap_3 PHY_8139 ();
 sky130_fd_sc_hd__decap_3 PHY_8140 ();
 sky130_fd_sc_hd__decap_3 PHY_8141 ();
 sky130_fd_sc_hd__decap_3 PHY_8142 ();
 sky130_fd_sc_hd__decap_3 PHY_8143 ();
 sky130_fd_sc_hd__decap_3 PHY_8144 ();
 sky130_fd_sc_hd__decap_3 PHY_8145 ();
 sky130_fd_sc_hd__decap_3 PHY_8146 ();
 sky130_fd_sc_hd__decap_3 PHY_8147 ();
 sky130_fd_sc_hd__decap_3 PHY_8148 ();
 sky130_fd_sc_hd__decap_3 PHY_8149 ();
 sky130_fd_sc_hd__decap_3 PHY_8150 ();
 sky130_fd_sc_hd__decap_3 PHY_8151 ();
 sky130_fd_sc_hd__decap_3 PHY_8152 ();
 sky130_fd_sc_hd__decap_3 PHY_8153 ();
 sky130_fd_sc_hd__decap_3 PHY_8154 ();
 sky130_fd_sc_hd__decap_3 PHY_8155 ();
 sky130_fd_sc_hd__decap_3 PHY_8156 ();
 sky130_fd_sc_hd__decap_3 PHY_8157 ();
 sky130_fd_sc_hd__decap_3 PHY_8158 ();
 sky130_fd_sc_hd__decap_3 PHY_8159 ();
 sky130_fd_sc_hd__decap_3 PHY_8160 ();
 sky130_fd_sc_hd__decap_3 PHY_8161 ();
 sky130_fd_sc_hd__decap_3 PHY_8162 ();
 sky130_fd_sc_hd__decap_3 PHY_8163 ();
 sky130_fd_sc_hd__decap_3 PHY_8164 ();
 sky130_fd_sc_hd__decap_3 PHY_8165 ();
 sky130_fd_sc_hd__decap_3 PHY_8166 ();
 sky130_fd_sc_hd__decap_3 PHY_8167 ();
 sky130_fd_sc_hd__decap_3 PHY_8168 ();
 sky130_fd_sc_hd__decap_3 PHY_8169 ();
 sky130_fd_sc_hd__decap_3 PHY_8170 ();
 sky130_fd_sc_hd__decap_3 PHY_8171 ();
 sky130_fd_sc_hd__decap_3 PHY_8172 ();
 sky130_fd_sc_hd__decap_3 PHY_8173 ();
 sky130_fd_sc_hd__decap_3 PHY_8174 ();
 sky130_fd_sc_hd__decap_3 PHY_8175 ();
 sky130_fd_sc_hd__decap_3 PHY_8176 ();
 sky130_fd_sc_hd__decap_3 PHY_8177 ();
 sky130_fd_sc_hd__decap_3 PHY_8178 ();
 sky130_fd_sc_hd__decap_3 PHY_8179 ();
 sky130_fd_sc_hd__decap_3 PHY_8180 ();
 sky130_fd_sc_hd__decap_3 PHY_8181 ();
 sky130_fd_sc_hd__decap_3 PHY_8182 ();
 sky130_fd_sc_hd__decap_3 PHY_8183 ();
 sky130_fd_sc_hd__decap_3 PHY_8184 ();
 sky130_fd_sc_hd__decap_3 PHY_8185 ();
 sky130_fd_sc_hd__decap_3 PHY_8186 ();
 sky130_fd_sc_hd__decap_3 PHY_8187 ();
 sky130_fd_sc_hd__decap_3 PHY_8188 ();
 sky130_fd_sc_hd__decap_3 PHY_8189 ();
 sky130_fd_sc_hd__decap_3 PHY_8190 ();
 sky130_fd_sc_hd__decap_3 PHY_8191 ();
 sky130_fd_sc_hd__decap_3 PHY_8192 ();
 sky130_fd_sc_hd__decap_3 PHY_8193 ();
 sky130_fd_sc_hd__decap_3 PHY_8194 ();
 sky130_fd_sc_hd__decap_3 PHY_8195 ();
 sky130_fd_sc_hd__decap_3 PHY_8196 ();
 sky130_fd_sc_hd__decap_3 PHY_8197 ();
 sky130_fd_sc_hd__decap_3 PHY_8198 ();
 sky130_fd_sc_hd__decap_3 PHY_8199 ();
 sky130_fd_sc_hd__decap_3 PHY_8200 ();
 sky130_fd_sc_hd__decap_3 PHY_8201 ();
 sky130_fd_sc_hd__decap_3 PHY_8202 ();
 sky130_fd_sc_hd__decap_3 PHY_8203 ();
 sky130_fd_sc_hd__decap_3 PHY_8204 ();
 sky130_fd_sc_hd__decap_3 PHY_8205 ();
 sky130_fd_sc_hd__decap_3 PHY_8206 ();
 sky130_fd_sc_hd__decap_3 PHY_8207 ();
 sky130_fd_sc_hd__decap_3 PHY_8208 ();
 sky130_fd_sc_hd__decap_3 PHY_8209 ();
 sky130_fd_sc_hd__decap_3 PHY_8210 ();
 sky130_fd_sc_hd__decap_3 PHY_8211 ();
 sky130_fd_sc_hd__decap_3 PHY_8212 ();
 sky130_fd_sc_hd__decap_3 PHY_8213 ();
 sky130_fd_sc_hd__decap_3 PHY_8214 ();
 sky130_fd_sc_hd__decap_3 PHY_8215 ();
 sky130_fd_sc_hd__decap_3 PHY_8216 ();
 sky130_fd_sc_hd__decap_3 PHY_8217 ();
 sky130_fd_sc_hd__decap_3 PHY_8218 ();
 sky130_fd_sc_hd__decap_3 PHY_8219 ();
 sky130_fd_sc_hd__decap_3 PHY_8220 ();
 sky130_fd_sc_hd__decap_3 PHY_8221 ();
 sky130_fd_sc_hd__decap_3 PHY_8222 ();
 sky130_fd_sc_hd__decap_3 PHY_8223 ();
 sky130_fd_sc_hd__decap_3 PHY_8224 ();
 sky130_fd_sc_hd__decap_3 PHY_8225 ();
 sky130_fd_sc_hd__decap_3 PHY_8226 ();
 sky130_fd_sc_hd__decap_3 PHY_8227 ();
 sky130_fd_sc_hd__decap_3 PHY_8228 ();
 sky130_fd_sc_hd__decap_3 PHY_8229 ();
 sky130_fd_sc_hd__decap_3 PHY_8230 ();
 sky130_fd_sc_hd__decap_3 PHY_8231 ();
 sky130_fd_sc_hd__decap_3 PHY_8232 ();
 sky130_fd_sc_hd__decap_3 PHY_8233 ();
 sky130_fd_sc_hd__decap_3 PHY_8234 ();
 sky130_fd_sc_hd__decap_3 PHY_8235 ();
 sky130_fd_sc_hd__decap_3 PHY_8236 ();
 sky130_fd_sc_hd__decap_3 PHY_8237 ();
 sky130_fd_sc_hd__decap_3 PHY_8238 ();
 sky130_fd_sc_hd__decap_3 PHY_8239 ();
 sky130_fd_sc_hd__decap_3 PHY_8240 ();
 sky130_fd_sc_hd__decap_3 PHY_8241 ();
 sky130_fd_sc_hd__decap_3 PHY_8242 ();
 sky130_fd_sc_hd__decap_3 PHY_8243 ();
 sky130_fd_sc_hd__decap_3 PHY_8244 ();
 sky130_fd_sc_hd__decap_3 PHY_8245 ();
 sky130_fd_sc_hd__decap_3 PHY_8246 ();
 sky130_fd_sc_hd__decap_3 PHY_8247 ();
 sky130_fd_sc_hd__decap_3 PHY_8248 ();
 sky130_fd_sc_hd__decap_3 PHY_8249 ();
 sky130_fd_sc_hd__decap_3 PHY_8250 ();
 sky130_fd_sc_hd__decap_3 PHY_8251 ();
 sky130_fd_sc_hd__decap_3 PHY_8252 ();
 sky130_fd_sc_hd__decap_3 PHY_8253 ();
 sky130_fd_sc_hd__decap_3 PHY_8254 ();
 sky130_fd_sc_hd__decap_3 PHY_8255 ();
 sky130_fd_sc_hd__decap_3 PHY_8256 ();
 sky130_fd_sc_hd__decap_3 PHY_8257 ();
 sky130_fd_sc_hd__decap_3 PHY_8258 ();
 sky130_fd_sc_hd__decap_3 PHY_8259 ();
 sky130_fd_sc_hd__decap_3 PHY_8260 ();
 sky130_fd_sc_hd__decap_3 PHY_8261 ();
 sky130_fd_sc_hd__decap_3 PHY_8262 ();
 sky130_fd_sc_hd__decap_3 PHY_8263 ();
 sky130_fd_sc_hd__decap_3 PHY_8264 ();
 sky130_fd_sc_hd__decap_3 PHY_8265 ();
 sky130_fd_sc_hd__decap_3 PHY_8266 ();
 sky130_fd_sc_hd__decap_3 PHY_8267 ();
 sky130_fd_sc_hd__decap_3 PHY_8268 ();
 sky130_fd_sc_hd__decap_3 PHY_8269 ();
 sky130_fd_sc_hd__decap_3 PHY_8270 ();
 sky130_fd_sc_hd__decap_3 PHY_8271 ();
 sky130_fd_sc_hd__decap_3 PHY_8272 ();
 sky130_fd_sc_hd__decap_3 PHY_8273 ();
 sky130_fd_sc_hd__decap_3 PHY_8274 ();
 sky130_fd_sc_hd__decap_3 PHY_8275 ();
 sky130_fd_sc_hd__decap_3 PHY_8276 ();
 sky130_fd_sc_hd__decap_3 PHY_8277 ();
 sky130_fd_sc_hd__decap_3 PHY_8278 ();
 sky130_fd_sc_hd__decap_3 PHY_8279 ();
 sky130_fd_sc_hd__decap_3 PHY_8280 ();
 sky130_fd_sc_hd__decap_3 PHY_8281 ();
 sky130_fd_sc_hd__decap_3 PHY_8282 ();
 sky130_fd_sc_hd__decap_3 PHY_8283 ();
 sky130_fd_sc_hd__decap_3 PHY_8284 ();
 sky130_fd_sc_hd__decap_3 PHY_8285 ();
 sky130_fd_sc_hd__decap_3 PHY_8286 ();
 sky130_fd_sc_hd__decap_3 PHY_8287 ();
 sky130_fd_sc_hd__decap_3 PHY_8288 ();
 sky130_fd_sc_hd__decap_3 PHY_8289 ();
 sky130_fd_sc_hd__decap_3 PHY_8290 ();
 sky130_fd_sc_hd__decap_3 PHY_8291 ();
 sky130_fd_sc_hd__decap_3 PHY_8292 ();
 sky130_fd_sc_hd__decap_3 PHY_8293 ();
 sky130_fd_sc_hd__decap_3 PHY_8294 ();
 sky130_fd_sc_hd__decap_3 PHY_8295 ();
 sky130_fd_sc_hd__decap_3 PHY_8296 ();
 sky130_fd_sc_hd__decap_3 PHY_8297 ();
 sky130_fd_sc_hd__decap_3 PHY_8298 ();
 sky130_fd_sc_hd__decap_3 PHY_8299 ();
 sky130_fd_sc_hd__decap_3 PHY_8300 ();
 sky130_fd_sc_hd__decap_3 PHY_8301 ();
 sky130_fd_sc_hd__decap_3 PHY_8302 ();
 sky130_fd_sc_hd__decap_3 PHY_8303 ();
 sky130_fd_sc_hd__decap_3 PHY_8304 ();
 sky130_fd_sc_hd__decap_3 PHY_8305 ();
 sky130_fd_sc_hd__decap_3 PHY_8306 ();
 sky130_fd_sc_hd__decap_3 PHY_8307 ();
 sky130_fd_sc_hd__decap_3 PHY_8308 ();
 sky130_fd_sc_hd__decap_3 PHY_8309 ();
 sky130_fd_sc_hd__decap_3 PHY_8310 ();
 sky130_fd_sc_hd__decap_3 PHY_8311 ();
 sky130_fd_sc_hd__decap_3 PHY_8312 ();
 sky130_fd_sc_hd__decap_3 PHY_8313 ();
 sky130_fd_sc_hd__decap_3 PHY_8314 ();
 sky130_fd_sc_hd__decap_3 PHY_8315 ();
 sky130_fd_sc_hd__decap_3 PHY_8316 ();
 sky130_fd_sc_hd__decap_3 PHY_8317 ();
 sky130_fd_sc_hd__decap_3 PHY_8318 ();
 sky130_fd_sc_hd__decap_3 PHY_8319 ();
 sky130_fd_sc_hd__decap_3 PHY_8320 ();
 sky130_fd_sc_hd__decap_3 PHY_8321 ();
 sky130_fd_sc_hd__decap_3 PHY_8322 ();
 sky130_fd_sc_hd__decap_3 PHY_8323 ();
 sky130_fd_sc_hd__decap_3 PHY_8324 ();
 sky130_fd_sc_hd__decap_3 PHY_8325 ();
 sky130_fd_sc_hd__decap_3 PHY_8326 ();
 sky130_fd_sc_hd__decap_3 PHY_8327 ();
 sky130_fd_sc_hd__decap_3 PHY_8328 ();
 sky130_fd_sc_hd__decap_3 PHY_8329 ();
 sky130_fd_sc_hd__decap_3 PHY_8330 ();
 sky130_fd_sc_hd__decap_3 PHY_8331 ();
 sky130_fd_sc_hd__decap_3 PHY_8332 ();
 sky130_fd_sc_hd__decap_3 PHY_8333 ();
 sky130_fd_sc_hd__decap_3 PHY_8334 ();
 sky130_fd_sc_hd__decap_3 PHY_8335 ();
 sky130_fd_sc_hd__decap_3 PHY_8336 ();
 sky130_fd_sc_hd__decap_3 PHY_8337 ();
 sky130_fd_sc_hd__decap_3 PHY_8338 ();
 sky130_fd_sc_hd__decap_3 PHY_8339 ();
 sky130_fd_sc_hd__decap_3 PHY_8340 ();
 sky130_fd_sc_hd__decap_3 PHY_8341 ();
 sky130_fd_sc_hd__decap_3 PHY_8342 ();
 sky130_fd_sc_hd__decap_3 PHY_8343 ();
 sky130_fd_sc_hd__decap_3 PHY_8344 ();
 sky130_fd_sc_hd__decap_3 PHY_8345 ();
 sky130_fd_sc_hd__decap_3 PHY_8346 ();
 sky130_fd_sc_hd__decap_3 PHY_8347 ();
 sky130_fd_sc_hd__decap_3 PHY_8348 ();
 sky130_fd_sc_hd__decap_3 PHY_8349 ();
 sky130_fd_sc_hd__decap_3 PHY_8350 ();
 sky130_fd_sc_hd__decap_3 PHY_8351 ();
 sky130_fd_sc_hd__decap_3 PHY_8352 ();
 sky130_fd_sc_hd__decap_3 PHY_8353 ();
 sky130_fd_sc_hd__decap_3 PHY_8354 ();
 sky130_fd_sc_hd__decap_3 PHY_8355 ();
 sky130_fd_sc_hd__decap_3 PHY_8356 ();
 sky130_fd_sc_hd__decap_3 PHY_8357 ();
 sky130_fd_sc_hd__decap_3 PHY_8358 ();
 sky130_fd_sc_hd__decap_3 PHY_8359 ();
 sky130_fd_sc_hd__decap_3 PHY_8360 ();
 sky130_fd_sc_hd__decap_3 PHY_8361 ();
 sky130_fd_sc_hd__decap_3 PHY_8362 ();
 sky130_fd_sc_hd__decap_3 PHY_8363 ();
 sky130_fd_sc_hd__decap_3 PHY_8364 ();
 sky130_fd_sc_hd__decap_3 PHY_8365 ();
 sky130_fd_sc_hd__decap_3 PHY_8366 ();
 sky130_fd_sc_hd__decap_3 PHY_8367 ();
 sky130_fd_sc_hd__decap_3 PHY_8368 ();
 sky130_fd_sc_hd__decap_3 PHY_8369 ();
 sky130_fd_sc_hd__decap_3 PHY_8370 ();
 sky130_fd_sc_hd__decap_3 PHY_8371 ();
 sky130_fd_sc_hd__decap_3 PHY_8372 ();
 sky130_fd_sc_hd__decap_3 PHY_8373 ();
 sky130_fd_sc_hd__decap_3 PHY_8374 ();
 sky130_fd_sc_hd__decap_3 PHY_8375 ();
 sky130_fd_sc_hd__decap_3 PHY_8376 ();
 sky130_fd_sc_hd__decap_3 PHY_8377 ();
 sky130_fd_sc_hd__decap_3 PHY_8378 ();
 sky130_fd_sc_hd__decap_3 PHY_8379 ();
 sky130_fd_sc_hd__decap_3 PHY_8380 ();
 sky130_fd_sc_hd__decap_3 PHY_8381 ();
 sky130_fd_sc_hd__decap_3 PHY_8382 ();
 sky130_fd_sc_hd__decap_3 PHY_8383 ();
 sky130_fd_sc_hd__decap_3 PHY_8384 ();
 sky130_fd_sc_hd__decap_3 PHY_8385 ();
 sky130_fd_sc_hd__decap_3 PHY_8386 ();
 sky130_fd_sc_hd__decap_3 PHY_8387 ();
 sky130_fd_sc_hd__decap_3 PHY_8388 ();
 sky130_fd_sc_hd__decap_3 PHY_8389 ();
 sky130_fd_sc_hd__decap_3 PHY_8390 ();
 sky130_fd_sc_hd__decap_3 PHY_8391 ();
 sky130_fd_sc_hd__decap_3 PHY_8392 ();
 sky130_fd_sc_hd__decap_3 PHY_8393 ();
 sky130_fd_sc_hd__decap_3 PHY_8394 ();
 sky130_fd_sc_hd__decap_3 PHY_8395 ();
 sky130_fd_sc_hd__decap_3 PHY_8396 ();
 sky130_fd_sc_hd__decap_3 PHY_8397 ();
 sky130_fd_sc_hd__decap_3 PHY_8398 ();
 sky130_fd_sc_hd__decap_3 PHY_8399 ();
 sky130_fd_sc_hd__decap_3 PHY_8400 ();
 sky130_fd_sc_hd__decap_3 PHY_8401 ();
 sky130_fd_sc_hd__decap_3 PHY_8402 ();
 sky130_fd_sc_hd__decap_3 PHY_8403 ();
 sky130_fd_sc_hd__decap_3 PHY_8404 ();
 sky130_fd_sc_hd__decap_3 PHY_8405 ();
 sky130_fd_sc_hd__decap_3 PHY_8406 ();
 sky130_fd_sc_hd__decap_3 PHY_8407 ();
 sky130_fd_sc_hd__decap_3 PHY_8408 ();
 sky130_fd_sc_hd__decap_3 PHY_8409 ();
 sky130_fd_sc_hd__decap_3 PHY_8410 ();
 sky130_fd_sc_hd__decap_3 PHY_8411 ();
 sky130_fd_sc_hd__decap_3 PHY_8412 ();
 sky130_fd_sc_hd__decap_3 PHY_8413 ();
 sky130_fd_sc_hd__decap_3 PHY_8414 ();
 sky130_fd_sc_hd__decap_3 PHY_8415 ();
 sky130_fd_sc_hd__decap_3 PHY_8416 ();
 sky130_fd_sc_hd__decap_3 PHY_8417 ();
 sky130_fd_sc_hd__decap_3 PHY_8418 ();
 sky130_fd_sc_hd__decap_3 PHY_8419 ();
 sky130_fd_sc_hd__decap_3 PHY_8420 ();
 sky130_fd_sc_hd__decap_3 PHY_8421 ();
 sky130_fd_sc_hd__decap_3 PHY_8422 ();
 sky130_fd_sc_hd__decap_3 PHY_8423 ();
 sky130_fd_sc_hd__decap_3 PHY_8424 ();
 sky130_fd_sc_hd__decap_3 PHY_8425 ();
 sky130_fd_sc_hd__decap_3 PHY_8426 ();
 sky130_fd_sc_hd__decap_3 PHY_8427 ();
 sky130_fd_sc_hd__decap_3 PHY_8428 ();
 sky130_fd_sc_hd__decap_3 PHY_8429 ();
 sky130_fd_sc_hd__decap_3 PHY_8430 ();
 sky130_fd_sc_hd__decap_3 PHY_8431 ();
 sky130_fd_sc_hd__decap_3 PHY_8432 ();
 sky130_fd_sc_hd__decap_3 PHY_8433 ();
 sky130_fd_sc_hd__decap_3 PHY_8434 ();
 sky130_fd_sc_hd__decap_3 PHY_8435 ();
 sky130_fd_sc_hd__decap_3 PHY_8436 ();
 sky130_fd_sc_hd__decap_3 PHY_8437 ();
 sky130_fd_sc_hd__decap_3 PHY_8438 ();
 sky130_fd_sc_hd__decap_3 PHY_8439 ();
 sky130_fd_sc_hd__decap_3 PHY_8440 ();
 sky130_fd_sc_hd__decap_3 PHY_8441 ();
 sky130_fd_sc_hd__decap_3 PHY_8442 ();
 sky130_fd_sc_hd__decap_3 PHY_8443 ();
 sky130_fd_sc_hd__decap_3 PHY_8444 ();
 sky130_fd_sc_hd__decap_3 PHY_8445 ();
 sky130_fd_sc_hd__decap_3 PHY_8446 ();
 sky130_fd_sc_hd__decap_3 PHY_8447 ();
 sky130_fd_sc_hd__decap_3 PHY_8448 ();
 sky130_fd_sc_hd__decap_3 PHY_8449 ();
 sky130_fd_sc_hd__decap_3 PHY_8450 ();
 sky130_fd_sc_hd__decap_3 PHY_8451 ();
 sky130_fd_sc_hd__decap_3 PHY_8452 ();
 sky130_fd_sc_hd__decap_3 PHY_8453 ();
 sky130_fd_sc_hd__decap_3 PHY_8454 ();
 sky130_fd_sc_hd__decap_3 PHY_8455 ();
 sky130_fd_sc_hd__decap_3 PHY_8456 ();
 sky130_fd_sc_hd__decap_3 PHY_8457 ();
 sky130_fd_sc_hd__decap_3 PHY_8458 ();
 sky130_fd_sc_hd__decap_3 PHY_8459 ();
 sky130_fd_sc_hd__decap_3 PHY_8460 ();
 sky130_fd_sc_hd__decap_3 PHY_8461 ();
 sky130_fd_sc_hd__decap_3 PHY_8462 ();
 sky130_fd_sc_hd__decap_3 PHY_8463 ();
 sky130_fd_sc_hd__decap_3 PHY_8464 ();
 sky130_fd_sc_hd__decap_3 PHY_8465 ();
 sky130_fd_sc_hd__decap_3 PHY_8466 ();
 sky130_fd_sc_hd__decap_3 PHY_8467 ();
 sky130_fd_sc_hd__decap_3 PHY_8468 ();
 sky130_fd_sc_hd__decap_3 PHY_8469 ();
 sky130_fd_sc_hd__decap_3 PHY_8470 ();
 sky130_fd_sc_hd__decap_3 PHY_8471 ();
 sky130_fd_sc_hd__decap_3 PHY_8472 ();
 sky130_fd_sc_hd__decap_3 PHY_8473 ();
 sky130_fd_sc_hd__decap_3 PHY_8474 ();
 sky130_fd_sc_hd__decap_3 PHY_8475 ();
 sky130_fd_sc_hd__decap_3 PHY_8476 ();
 sky130_fd_sc_hd__decap_3 PHY_8477 ();
 sky130_fd_sc_hd__decap_3 PHY_8478 ();
 sky130_fd_sc_hd__decap_3 PHY_8479 ();
 sky130_fd_sc_hd__decap_3 PHY_8480 ();
 sky130_fd_sc_hd__decap_3 PHY_8481 ();
 sky130_fd_sc_hd__decap_3 PHY_8482 ();
 sky130_fd_sc_hd__decap_3 PHY_8483 ();
 sky130_fd_sc_hd__decap_3 PHY_8484 ();
 sky130_fd_sc_hd__decap_3 PHY_8485 ();
 sky130_fd_sc_hd__decap_3 PHY_8486 ();
 sky130_fd_sc_hd__decap_3 PHY_8487 ();
 sky130_fd_sc_hd__decap_3 PHY_8488 ();
 sky130_fd_sc_hd__decap_3 PHY_8489 ();
 sky130_fd_sc_hd__decap_3 PHY_8490 ();
 sky130_fd_sc_hd__decap_3 PHY_8491 ();
 sky130_fd_sc_hd__decap_3 PHY_8492 ();
 sky130_fd_sc_hd__decap_3 PHY_8493 ();
 sky130_fd_sc_hd__decap_3 PHY_8494 ();
 sky130_fd_sc_hd__decap_3 PHY_8495 ();
 sky130_fd_sc_hd__decap_3 PHY_8496 ();
 sky130_fd_sc_hd__decap_3 PHY_8497 ();
 sky130_fd_sc_hd__decap_3 PHY_8498 ();
 sky130_fd_sc_hd__decap_3 PHY_8499 ();
 sky130_fd_sc_hd__decap_3 PHY_8500 ();
 sky130_fd_sc_hd__decap_3 PHY_8501 ();
 sky130_fd_sc_hd__decap_3 PHY_8502 ();
 sky130_fd_sc_hd__decap_3 PHY_8503 ();
 sky130_fd_sc_hd__decap_3 PHY_8504 ();
 sky130_fd_sc_hd__decap_3 PHY_8505 ();
 sky130_fd_sc_hd__decap_3 PHY_8506 ();
 sky130_fd_sc_hd__decap_3 PHY_8507 ();
 sky130_fd_sc_hd__decap_3 PHY_8508 ();
 sky130_fd_sc_hd__decap_3 PHY_8509 ();
 sky130_fd_sc_hd__decap_3 PHY_8510 ();
 sky130_fd_sc_hd__decap_3 PHY_8511 ();
 sky130_fd_sc_hd__decap_3 PHY_8512 ();
 sky130_fd_sc_hd__decap_3 PHY_8513 ();
 sky130_fd_sc_hd__decap_3 PHY_8514 ();
 sky130_fd_sc_hd__decap_3 PHY_8515 ();
 sky130_fd_sc_hd__decap_3 PHY_8516 ();
 sky130_fd_sc_hd__decap_3 PHY_8517 ();
 sky130_fd_sc_hd__decap_3 PHY_8518 ();
 sky130_fd_sc_hd__decap_3 PHY_8519 ();
 sky130_fd_sc_hd__decap_3 PHY_8520 ();
 sky130_fd_sc_hd__decap_3 PHY_8521 ();
 sky130_fd_sc_hd__decap_3 PHY_8522 ();
 sky130_fd_sc_hd__decap_3 PHY_8523 ();
 sky130_fd_sc_hd__decap_3 PHY_8524 ();
 sky130_fd_sc_hd__decap_3 PHY_8525 ();
 sky130_fd_sc_hd__decap_3 PHY_8526 ();
 sky130_fd_sc_hd__decap_3 PHY_8527 ();
 sky130_fd_sc_hd__decap_3 PHY_8528 ();
 sky130_fd_sc_hd__decap_3 PHY_8529 ();
 sky130_fd_sc_hd__decap_3 PHY_8530 ();
 sky130_fd_sc_hd__decap_3 PHY_8531 ();
 sky130_fd_sc_hd__decap_3 PHY_8532 ();
 sky130_fd_sc_hd__decap_3 PHY_8533 ();
 sky130_fd_sc_hd__decap_3 PHY_8534 ();
 sky130_fd_sc_hd__decap_3 PHY_8535 ();
 sky130_fd_sc_hd__decap_3 PHY_8536 ();
 sky130_fd_sc_hd__decap_3 PHY_8537 ();
 sky130_fd_sc_hd__decap_3 PHY_8538 ();
 sky130_fd_sc_hd__decap_3 PHY_8539 ();
 sky130_fd_sc_hd__decap_3 PHY_8540 ();
 sky130_fd_sc_hd__decap_3 PHY_8541 ();
 sky130_fd_sc_hd__decap_3 PHY_8542 ();
 sky130_fd_sc_hd__decap_3 PHY_8543 ();
 sky130_fd_sc_hd__decap_3 PHY_8544 ();
 sky130_fd_sc_hd__decap_3 PHY_8545 ();
 sky130_fd_sc_hd__decap_3 PHY_8546 ();
 sky130_fd_sc_hd__decap_3 PHY_8547 ();
 sky130_fd_sc_hd__decap_3 PHY_8548 ();
 sky130_fd_sc_hd__decap_3 PHY_8549 ();
 sky130_fd_sc_hd__decap_3 PHY_8550 ();
 sky130_fd_sc_hd__decap_3 PHY_8551 ();
 sky130_fd_sc_hd__decap_3 PHY_8552 ();
 sky130_fd_sc_hd__decap_3 PHY_8553 ();
 sky130_fd_sc_hd__decap_3 PHY_8554 ();
 sky130_fd_sc_hd__decap_3 PHY_8555 ();
 sky130_fd_sc_hd__decap_3 PHY_8556 ();
 sky130_fd_sc_hd__decap_3 PHY_8557 ();
 sky130_fd_sc_hd__decap_3 PHY_8558 ();
 sky130_fd_sc_hd__decap_3 PHY_8559 ();
 sky130_fd_sc_hd__decap_3 PHY_8560 ();
 sky130_fd_sc_hd__decap_3 PHY_8561 ();
 sky130_fd_sc_hd__decap_3 PHY_8562 ();
 sky130_fd_sc_hd__decap_3 PHY_8563 ();
 sky130_fd_sc_hd__decap_3 PHY_8564 ();
 sky130_fd_sc_hd__decap_3 PHY_8565 ();
 sky130_fd_sc_hd__decap_3 PHY_8566 ();
 sky130_fd_sc_hd__decap_3 PHY_8567 ();
 sky130_fd_sc_hd__decap_3 PHY_8568 ();
 sky130_fd_sc_hd__decap_3 PHY_8569 ();
 sky130_fd_sc_hd__decap_3 PHY_8570 ();
 sky130_fd_sc_hd__decap_3 PHY_8571 ();
 sky130_fd_sc_hd__decap_3 PHY_8572 ();
 sky130_fd_sc_hd__decap_3 PHY_8573 ();
 sky130_fd_sc_hd__decap_3 PHY_8574 ();
 sky130_fd_sc_hd__decap_3 PHY_8575 ();
 sky130_fd_sc_hd__decap_3 PHY_8576 ();
 sky130_fd_sc_hd__decap_3 PHY_8577 ();
 sky130_fd_sc_hd__decap_3 PHY_8578 ();
 sky130_fd_sc_hd__decap_3 PHY_8579 ();
 sky130_fd_sc_hd__decap_3 PHY_8580 ();
 sky130_fd_sc_hd__decap_3 PHY_8581 ();
 sky130_fd_sc_hd__decap_3 PHY_8582 ();
 sky130_fd_sc_hd__decap_3 PHY_8583 ();
 sky130_fd_sc_hd__decap_3 PHY_8584 ();
 sky130_fd_sc_hd__decap_3 PHY_8585 ();
 sky130_fd_sc_hd__decap_3 PHY_8586 ();
 sky130_fd_sc_hd__decap_3 PHY_8587 ();
 sky130_fd_sc_hd__decap_3 PHY_8588 ();
 sky130_fd_sc_hd__decap_3 PHY_8589 ();
 sky130_fd_sc_hd__decap_3 PHY_8590 ();
 sky130_fd_sc_hd__decap_3 PHY_8591 ();
 sky130_fd_sc_hd__decap_3 PHY_8592 ();
 sky130_fd_sc_hd__decap_3 PHY_8593 ();
 sky130_fd_sc_hd__decap_3 PHY_8594 ();
 sky130_fd_sc_hd__decap_3 PHY_8595 ();
 sky130_fd_sc_hd__decap_3 PHY_8596 ();
 sky130_fd_sc_hd__decap_3 PHY_8597 ();
 sky130_fd_sc_hd__decap_3 PHY_8598 ();
 sky130_fd_sc_hd__decap_3 PHY_8599 ();
 sky130_fd_sc_hd__decap_3 PHY_8600 ();
 sky130_fd_sc_hd__decap_3 PHY_8601 ();
 sky130_fd_sc_hd__decap_3 PHY_8602 ();
 sky130_fd_sc_hd__decap_3 PHY_8603 ();
 sky130_fd_sc_hd__decap_3 PHY_8604 ();
 sky130_fd_sc_hd__decap_3 PHY_8605 ();
 sky130_fd_sc_hd__decap_3 PHY_8606 ();
 sky130_fd_sc_hd__decap_3 PHY_8607 ();
 sky130_fd_sc_hd__decap_3 PHY_8608 ();
 sky130_fd_sc_hd__decap_3 PHY_8609 ();
 sky130_fd_sc_hd__decap_3 PHY_8610 ();
 sky130_fd_sc_hd__decap_3 PHY_8611 ();
 sky130_fd_sc_hd__decap_3 PHY_8612 ();
 sky130_fd_sc_hd__decap_3 PHY_8613 ();
 sky130_fd_sc_hd__decap_3 PHY_8614 ();
 sky130_fd_sc_hd__decap_3 PHY_8615 ();
 sky130_fd_sc_hd__decap_3 PHY_8616 ();
 sky130_fd_sc_hd__decap_3 PHY_8617 ();
 sky130_fd_sc_hd__decap_3 PHY_8618 ();
 sky130_fd_sc_hd__decap_3 PHY_8619 ();
 sky130_fd_sc_hd__decap_3 PHY_8620 ();
 sky130_fd_sc_hd__decap_3 PHY_8621 ();
 sky130_fd_sc_hd__decap_3 PHY_8622 ();
 sky130_fd_sc_hd__decap_3 PHY_8623 ();
 sky130_fd_sc_hd__decap_3 PHY_8624 ();
 sky130_fd_sc_hd__decap_3 PHY_8625 ();
 sky130_fd_sc_hd__decap_3 PHY_8626 ();
 sky130_fd_sc_hd__decap_3 PHY_8627 ();
 sky130_fd_sc_hd__decap_3 PHY_8628 ();
 sky130_fd_sc_hd__decap_3 PHY_8629 ();
 sky130_fd_sc_hd__decap_3 PHY_8630 ();
 sky130_fd_sc_hd__decap_3 PHY_8631 ();
 sky130_fd_sc_hd__decap_3 PHY_8632 ();
 sky130_fd_sc_hd__decap_3 PHY_8633 ();
 sky130_fd_sc_hd__decap_3 PHY_8634 ();
 sky130_fd_sc_hd__decap_3 PHY_8635 ();
 sky130_fd_sc_hd__decap_3 PHY_8636 ();
 sky130_fd_sc_hd__decap_3 PHY_8637 ();
 sky130_fd_sc_hd__decap_3 PHY_8638 ();
 sky130_fd_sc_hd__decap_3 PHY_8639 ();
 sky130_fd_sc_hd__decap_3 PHY_8640 ();
 sky130_fd_sc_hd__decap_3 PHY_8641 ();
 sky130_fd_sc_hd__decap_3 PHY_8642 ();
 sky130_fd_sc_hd__decap_3 PHY_8643 ();
 sky130_fd_sc_hd__decap_3 PHY_8644 ();
 sky130_fd_sc_hd__decap_3 PHY_8645 ();
 sky130_fd_sc_hd__decap_3 PHY_8646 ();
 sky130_fd_sc_hd__decap_3 PHY_8647 ();
 sky130_fd_sc_hd__decap_3 PHY_8648 ();
 sky130_fd_sc_hd__decap_3 PHY_8649 ();
 sky130_fd_sc_hd__decap_3 PHY_8650 ();
 sky130_fd_sc_hd__decap_3 PHY_8651 ();
 sky130_fd_sc_hd__decap_3 PHY_8652 ();
 sky130_fd_sc_hd__decap_3 PHY_8653 ();
 sky130_fd_sc_hd__decap_3 PHY_8654 ();
 sky130_fd_sc_hd__decap_3 PHY_8655 ();
 sky130_fd_sc_hd__decap_3 PHY_8656 ();
 sky130_fd_sc_hd__decap_3 PHY_8657 ();
 sky130_fd_sc_hd__decap_3 PHY_8658 ();
 sky130_fd_sc_hd__decap_3 PHY_8659 ();
 sky130_fd_sc_hd__decap_3 PHY_8660 ();
 sky130_fd_sc_hd__decap_3 PHY_8661 ();
 sky130_fd_sc_hd__decap_3 PHY_8662 ();
 sky130_fd_sc_hd__decap_3 PHY_8663 ();
 sky130_fd_sc_hd__decap_3 PHY_8664 ();
 sky130_fd_sc_hd__decap_3 PHY_8665 ();
 sky130_fd_sc_hd__decap_3 PHY_8666 ();
 sky130_fd_sc_hd__decap_3 PHY_8667 ();
 sky130_fd_sc_hd__decap_3 PHY_8668 ();
 sky130_fd_sc_hd__decap_3 PHY_8669 ();
 sky130_fd_sc_hd__decap_3 PHY_8670 ();
 sky130_fd_sc_hd__decap_3 PHY_8671 ();
 sky130_fd_sc_hd__decap_3 PHY_8672 ();
 sky130_fd_sc_hd__decap_3 PHY_8673 ();
 sky130_fd_sc_hd__decap_3 PHY_8674 ();
 sky130_fd_sc_hd__decap_3 PHY_8675 ();
 sky130_fd_sc_hd__decap_3 PHY_8676 ();
 sky130_fd_sc_hd__decap_3 PHY_8677 ();
 sky130_fd_sc_hd__decap_3 PHY_8678 ();
 sky130_fd_sc_hd__decap_3 PHY_8679 ();
 sky130_fd_sc_hd__decap_3 PHY_8680 ();
 sky130_fd_sc_hd__decap_3 PHY_8681 ();
 sky130_fd_sc_hd__decap_3 PHY_8682 ();
 sky130_fd_sc_hd__decap_3 PHY_8683 ();
 sky130_fd_sc_hd__decap_3 PHY_8684 ();
 sky130_fd_sc_hd__decap_3 PHY_8685 ();
 sky130_fd_sc_hd__decap_3 PHY_8686 ();
 sky130_fd_sc_hd__decap_3 PHY_8687 ();
 sky130_fd_sc_hd__decap_3 PHY_8688 ();
 sky130_fd_sc_hd__decap_3 PHY_8689 ();
 sky130_fd_sc_hd__decap_3 PHY_8690 ();
 sky130_fd_sc_hd__decap_3 PHY_8691 ();
 sky130_fd_sc_hd__decap_3 PHY_8692 ();
 sky130_fd_sc_hd__decap_3 PHY_8693 ();
 sky130_fd_sc_hd__decap_3 PHY_8694 ();
 sky130_fd_sc_hd__decap_3 PHY_8695 ();
 sky130_fd_sc_hd__decap_3 PHY_8696 ();
 sky130_fd_sc_hd__decap_3 PHY_8697 ();
 sky130_fd_sc_hd__decap_3 PHY_8698 ();
 sky130_fd_sc_hd__decap_3 PHY_8699 ();
 sky130_fd_sc_hd__decap_3 PHY_8700 ();
 sky130_fd_sc_hd__decap_3 PHY_8701 ();
 sky130_fd_sc_hd__decap_3 PHY_8702 ();
 sky130_fd_sc_hd__decap_3 PHY_8703 ();
 sky130_fd_sc_hd__decap_3 PHY_8704 ();
 sky130_fd_sc_hd__decap_3 PHY_8705 ();
 sky130_fd_sc_hd__decap_3 PHY_8706 ();
 sky130_fd_sc_hd__decap_3 PHY_8707 ();
 sky130_fd_sc_hd__decap_3 PHY_8708 ();
 sky130_fd_sc_hd__decap_3 PHY_8709 ();
 sky130_fd_sc_hd__decap_3 PHY_8710 ();
 sky130_fd_sc_hd__decap_3 PHY_8711 ();
 sky130_fd_sc_hd__decap_3 PHY_8712 ();
 sky130_fd_sc_hd__decap_3 PHY_8713 ();
 sky130_fd_sc_hd__decap_3 PHY_8714 ();
 sky130_fd_sc_hd__decap_3 PHY_8715 ();
 sky130_fd_sc_hd__decap_3 PHY_8716 ();
 sky130_fd_sc_hd__decap_3 PHY_8717 ();
 sky130_fd_sc_hd__decap_3 PHY_8718 ();
 sky130_fd_sc_hd__decap_3 PHY_8719 ();
 sky130_fd_sc_hd__decap_3 PHY_8720 ();
 sky130_fd_sc_hd__decap_3 PHY_8721 ();
 sky130_fd_sc_hd__decap_3 PHY_8722 ();
 sky130_fd_sc_hd__decap_3 PHY_8723 ();
 sky130_fd_sc_hd__decap_3 PHY_8724 ();
 sky130_fd_sc_hd__decap_3 PHY_8725 ();
 sky130_fd_sc_hd__decap_3 PHY_8726 ();
 sky130_fd_sc_hd__decap_3 PHY_8727 ();
 sky130_fd_sc_hd__decap_3 PHY_8728 ();
 sky130_fd_sc_hd__decap_3 PHY_8729 ();
 sky130_fd_sc_hd__decap_3 PHY_8730 ();
 sky130_fd_sc_hd__decap_3 PHY_8731 ();
 sky130_fd_sc_hd__decap_3 PHY_8732 ();
 sky130_fd_sc_hd__decap_3 PHY_8733 ();
 sky130_fd_sc_hd__decap_3 PHY_8734 ();
 sky130_fd_sc_hd__decap_3 PHY_8735 ();
 sky130_fd_sc_hd__decap_3 PHY_8736 ();
 sky130_fd_sc_hd__decap_3 PHY_8737 ();
 sky130_fd_sc_hd__decap_3 PHY_8738 ();
 sky130_fd_sc_hd__decap_3 PHY_8739 ();
 sky130_fd_sc_hd__decap_3 PHY_8740 ();
 sky130_fd_sc_hd__decap_3 PHY_8741 ();
 sky130_fd_sc_hd__decap_3 PHY_8742 ();
 sky130_fd_sc_hd__decap_3 PHY_8743 ();
 sky130_fd_sc_hd__decap_3 PHY_8744 ();
 sky130_fd_sc_hd__decap_3 PHY_8745 ();
 sky130_fd_sc_hd__decap_3 PHY_8746 ();
 sky130_fd_sc_hd__decap_3 PHY_8747 ();
 sky130_fd_sc_hd__decap_3 PHY_8748 ();
 sky130_fd_sc_hd__decap_3 PHY_8749 ();
 sky130_fd_sc_hd__decap_3 PHY_8750 ();
 sky130_fd_sc_hd__decap_3 PHY_8751 ();
 sky130_fd_sc_hd__decap_3 PHY_8752 ();
 sky130_fd_sc_hd__decap_3 PHY_8753 ();
 sky130_fd_sc_hd__decap_3 PHY_8754 ();
 sky130_fd_sc_hd__decap_3 PHY_8755 ();
 sky130_fd_sc_hd__decap_3 PHY_8756 ();
 sky130_fd_sc_hd__decap_3 PHY_8757 ();
 sky130_fd_sc_hd__decap_3 PHY_8758 ();
 sky130_fd_sc_hd__decap_3 PHY_8759 ();
 sky130_fd_sc_hd__decap_3 PHY_8760 ();
 sky130_fd_sc_hd__decap_3 PHY_8761 ();
 sky130_fd_sc_hd__decap_3 PHY_8762 ();
 sky130_fd_sc_hd__decap_3 PHY_8763 ();
 sky130_fd_sc_hd__decap_3 PHY_8764 ();
 sky130_fd_sc_hd__decap_3 PHY_8765 ();
 sky130_fd_sc_hd__decap_3 PHY_8766 ();
 sky130_fd_sc_hd__decap_3 PHY_8767 ();
 sky130_fd_sc_hd__decap_3 PHY_8768 ();
 sky130_fd_sc_hd__decap_3 PHY_8769 ();
 sky130_fd_sc_hd__decap_3 PHY_8770 ();
 sky130_fd_sc_hd__decap_3 PHY_8771 ();
 sky130_fd_sc_hd__decap_3 PHY_8772 ();
 sky130_fd_sc_hd__decap_3 PHY_8773 ();
 sky130_fd_sc_hd__decap_3 PHY_8774 ();
 sky130_fd_sc_hd__decap_3 PHY_8775 ();
 sky130_fd_sc_hd__decap_3 PHY_8776 ();
 sky130_fd_sc_hd__decap_3 PHY_8777 ();
 sky130_fd_sc_hd__decap_3 PHY_8778 ();
 sky130_fd_sc_hd__decap_3 PHY_8779 ();
 sky130_fd_sc_hd__decap_3 PHY_8780 ();
 sky130_fd_sc_hd__decap_3 PHY_8781 ();
 sky130_fd_sc_hd__decap_3 PHY_8782 ();
 sky130_fd_sc_hd__decap_3 PHY_8783 ();
 sky130_fd_sc_hd__decap_3 PHY_8784 ();
 sky130_fd_sc_hd__decap_3 PHY_8785 ();
 sky130_fd_sc_hd__decap_3 PHY_8786 ();
 sky130_fd_sc_hd__decap_3 PHY_8787 ();
 sky130_fd_sc_hd__decap_3 PHY_8788 ();
 sky130_fd_sc_hd__decap_3 PHY_8789 ();
 sky130_fd_sc_hd__decap_3 PHY_8790 ();
 sky130_fd_sc_hd__decap_3 PHY_8791 ();
 sky130_fd_sc_hd__decap_3 PHY_8792 ();
 sky130_fd_sc_hd__decap_3 PHY_8793 ();
 sky130_fd_sc_hd__decap_3 PHY_8794 ();
 sky130_fd_sc_hd__decap_3 PHY_8795 ();
 sky130_fd_sc_hd__decap_3 PHY_8796 ();
 sky130_fd_sc_hd__decap_3 PHY_8797 ();
 sky130_fd_sc_hd__decap_3 PHY_8798 ();
 sky130_fd_sc_hd__decap_3 PHY_8799 ();
 sky130_fd_sc_hd__decap_3 PHY_8800 ();
 sky130_fd_sc_hd__decap_3 PHY_8801 ();
 sky130_fd_sc_hd__decap_3 PHY_8802 ();
 sky130_fd_sc_hd__decap_3 PHY_8803 ();
 sky130_fd_sc_hd__decap_3 PHY_8804 ();
 sky130_fd_sc_hd__decap_3 PHY_8805 ();
 sky130_fd_sc_hd__decap_3 PHY_8806 ();
 sky130_fd_sc_hd__decap_3 PHY_8807 ();
 sky130_fd_sc_hd__decap_3 PHY_8808 ();
 sky130_fd_sc_hd__decap_3 PHY_8809 ();
 sky130_fd_sc_hd__decap_3 PHY_8810 ();
 sky130_fd_sc_hd__decap_3 PHY_8811 ();
 sky130_fd_sc_hd__decap_3 PHY_8812 ();
 sky130_fd_sc_hd__decap_3 PHY_8813 ();
 sky130_fd_sc_hd__decap_3 PHY_8814 ();
 sky130_fd_sc_hd__decap_3 PHY_8815 ();
 sky130_fd_sc_hd__decap_3 PHY_8816 ();
 sky130_fd_sc_hd__decap_3 PHY_8817 ();
 sky130_fd_sc_hd__decap_3 PHY_8818 ();
 sky130_fd_sc_hd__decap_3 PHY_8819 ();
 sky130_fd_sc_hd__decap_3 PHY_8820 ();
 sky130_fd_sc_hd__decap_3 PHY_8821 ();
 sky130_fd_sc_hd__decap_3 PHY_8822 ();
 sky130_fd_sc_hd__decap_3 PHY_8823 ();
 sky130_fd_sc_hd__decap_3 PHY_8824 ();
 sky130_fd_sc_hd__decap_3 PHY_8825 ();
 sky130_fd_sc_hd__decap_3 PHY_8826 ();
 sky130_fd_sc_hd__decap_3 PHY_8827 ();
 sky130_fd_sc_hd__decap_3 PHY_8828 ();
 sky130_fd_sc_hd__decap_3 PHY_8829 ();
 sky130_fd_sc_hd__decap_3 PHY_8830 ();
 sky130_fd_sc_hd__decap_3 PHY_8831 ();
 sky130_fd_sc_hd__decap_3 PHY_8832 ();
 sky130_fd_sc_hd__decap_3 PHY_8833 ();
 sky130_fd_sc_hd__decap_3 PHY_8834 ();
 sky130_fd_sc_hd__decap_3 PHY_8835 ();
 sky130_fd_sc_hd__decap_3 PHY_8836 ();
 sky130_fd_sc_hd__decap_3 PHY_8837 ();
 sky130_fd_sc_hd__decap_3 PHY_8838 ();
 sky130_fd_sc_hd__decap_3 PHY_8839 ();
 sky130_fd_sc_hd__decap_3 PHY_8840 ();
 sky130_fd_sc_hd__decap_3 PHY_8841 ();
 sky130_fd_sc_hd__decap_3 PHY_8842 ();
 sky130_fd_sc_hd__decap_3 PHY_8843 ();
 sky130_fd_sc_hd__decap_3 PHY_8844 ();
 sky130_fd_sc_hd__decap_3 PHY_8845 ();
 sky130_fd_sc_hd__decap_3 PHY_8846 ();
 sky130_fd_sc_hd__decap_3 PHY_8847 ();
 sky130_fd_sc_hd__decap_3 PHY_8848 ();
 sky130_fd_sc_hd__decap_3 PHY_8849 ();
 sky130_fd_sc_hd__decap_3 PHY_8850 ();
 sky130_fd_sc_hd__decap_3 PHY_8851 ();
 sky130_fd_sc_hd__decap_3 PHY_8852 ();
 sky130_fd_sc_hd__decap_3 PHY_8853 ();
 sky130_fd_sc_hd__decap_3 PHY_8854 ();
 sky130_fd_sc_hd__decap_3 PHY_8855 ();
 sky130_fd_sc_hd__decap_3 PHY_8856 ();
 sky130_fd_sc_hd__decap_3 PHY_8857 ();
 sky130_fd_sc_hd__decap_3 PHY_8858 ();
 sky130_fd_sc_hd__decap_3 PHY_8859 ();
 sky130_fd_sc_hd__decap_3 PHY_8860 ();
 sky130_fd_sc_hd__decap_3 PHY_8861 ();
 sky130_fd_sc_hd__decap_3 PHY_8862 ();
 sky130_fd_sc_hd__decap_3 PHY_8863 ();
 sky130_fd_sc_hd__decap_3 PHY_8864 ();
 sky130_fd_sc_hd__decap_3 PHY_8865 ();
 sky130_fd_sc_hd__decap_3 PHY_8866 ();
 sky130_fd_sc_hd__decap_3 PHY_8867 ();
 sky130_fd_sc_hd__decap_3 PHY_8868 ();
 sky130_fd_sc_hd__decap_3 PHY_8869 ();
 sky130_fd_sc_hd__decap_3 PHY_8870 ();
 sky130_fd_sc_hd__decap_3 PHY_8871 ();
 sky130_fd_sc_hd__decap_3 PHY_8872 ();
 sky130_fd_sc_hd__decap_3 PHY_8873 ();
 sky130_fd_sc_hd__decap_3 PHY_8874 ();
 sky130_fd_sc_hd__decap_3 PHY_8875 ();
 sky130_fd_sc_hd__decap_3 PHY_8876 ();
 sky130_fd_sc_hd__decap_3 PHY_8877 ();
 sky130_fd_sc_hd__decap_3 PHY_8878 ();
 sky130_fd_sc_hd__decap_3 PHY_8879 ();
 sky130_fd_sc_hd__decap_3 PHY_8880 ();
 sky130_fd_sc_hd__decap_3 PHY_8881 ();
 sky130_fd_sc_hd__decap_3 PHY_8882 ();
 sky130_fd_sc_hd__decap_3 PHY_8883 ();
 sky130_fd_sc_hd__decap_3 PHY_8884 ();
 sky130_fd_sc_hd__decap_3 PHY_8885 ();
 sky130_fd_sc_hd__decap_3 PHY_8886 ();
 sky130_fd_sc_hd__decap_3 PHY_8887 ();
 sky130_fd_sc_hd__decap_3 PHY_8888 ();
 sky130_fd_sc_hd__decap_3 PHY_8889 ();
 sky130_fd_sc_hd__decap_3 PHY_8890 ();
 sky130_fd_sc_hd__decap_3 PHY_8891 ();
 sky130_fd_sc_hd__decap_3 PHY_8892 ();
 sky130_fd_sc_hd__decap_3 PHY_8893 ();
 sky130_fd_sc_hd__decap_3 PHY_8894 ();
 sky130_fd_sc_hd__decap_3 PHY_8895 ();
 sky130_fd_sc_hd__decap_3 PHY_8896 ();
 sky130_fd_sc_hd__decap_3 PHY_8897 ();
 sky130_fd_sc_hd__decap_3 PHY_8898 ();
 sky130_fd_sc_hd__decap_3 PHY_8899 ();
 sky130_fd_sc_hd__decap_3 PHY_8900 ();
 sky130_fd_sc_hd__decap_3 PHY_8901 ();
 sky130_fd_sc_hd__decap_3 PHY_8902 ();
 sky130_fd_sc_hd__decap_3 PHY_8903 ();
 sky130_fd_sc_hd__decap_3 PHY_8904 ();
 sky130_fd_sc_hd__decap_3 PHY_8905 ();
 sky130_fd_sc_hd__decap_3 PHY_8906 ();
 sky130_fd_sc_hd__decap_3 PHY_8907 ();
 sky130_fd_sc_hd__decap_3 PHY_8908 ();
 sky130_fd_sc_hd__decap_3 PHY_8909 ();
 sky130_fd_sc_hd__decap_3 PHY_8910 ();
 sky130_fd_sc_hd__decap_3 PHY_8911 ();
 sky130_fd_sc_hd__decap_3 PHY_8912 ();
 sky130_fd_sc_hd__decap_3 PHY_8913 ();
 sky130_fd_sc_hd__decap_3 PHY_8914 ();
 sky130_fd_sc_hd__decap_3 PHY_8915 ();
 sky130_fd_sc_hd__decap_3 PHY_8916 ();
 sky130_fd_sc_hd__decap_3 PHY_8917 ();
 sky130_fd_sc_hd__decap_3 PHY_8918 ();
 sky130_fd_sc_hd__decap_3 PHY_8919 ();
 sky130_fd_sc_hd__decap_3 PHY_8920 ();
 sky130_fd_sc_hd__decap_3 PHY_8921 ();
 sky130_fd_sc_hd__decap_3 PHY_8922 ();
 sky130_fd_sc_hd__decap_3 PHY_8923 ();
 sky130_fd_sc_hd__decap_3 PHY_8924 ();
 sky130_fd_sc_hd__decap_3 PHY_8925 ();
 sky130_fd_sc_hd__decap_3 PHY_8926 ();
 sky130_fd_sc_hd__decap_3 PHY_8927 ();
 sky130_fd_sc_hd__decap_3 PHY_8928 ();
 sky130_fd_sc_hd__decap_3 PHY_8929 ();
 sky130_fd_sc_hd__decap_3 PHY_8930 ();
 sky130_fd_sc_hd__decap_3 PHY_8931 ();
 sky130_fd_sc_hd__decap_3 PHY_8932 ();
 sky130_fd_sc_hd__decap_3 PHY_8933 ();
 sky130_fd_sc_hd__decap_3 PHY_8934 ();
 sky130_fd_sc_hd__decap_3 PHY_8935 ();
 sky130_fd_sc_hd__decap_3 PHY_8936 ();
 sky130_fd_sc_hd__decap_3 PHY_8937 ();
 sky130_fd_sc_hd__decap_3 PHY_8938 ();
 sky130_fd_sc_hd__decap_3 PHY_8939 ();
 sky130_fd_sc_hd__decap_3 PHY_8940 ();
 sky130_fd_sc_hd__decap_3 PHY_8941 ();
 sky130_fd_sc_hd__decap_3 PHY_8942 ();
 sky130_fd_sc_hd__decap_3 PHY_8943 ();
 sky130_fd_sc_hd__decap_3 PHY_8944 ();
 sky130_fd_sc_hd__decap_3 PHY_8945 ();
 sky130_fd_sc_hd__decap_3 PHY_8946 ();
 sky130_fd_sc_hd__decap_3 PHY_8947 ();
 sky130_fd_sc_hd__decap_3 PHY_8948 ();
 sky130_fd_sc_hd__decap_3 PHY_8949 ();
 sky130_fd_sc_hd__decap_3 PHY_8950 ();
 sky130_fd_sc_hd__decap_3 PHY_8951 ();
 sky130_fd_sc_hd__decap_3 PHY_8952 ();
 sky130_fd_sc_hd__decap_3 PHY_8953 ();
 sky130_fd_sc_hd__decap_3 PHY_8954 ();
 sky130_fd_sc_hd__decap_3 PHY_8955 ();
 sky130_fd_sc_hd__decap_3 PHY_8956 ();
 sky130_fd_sc_hd__decap_3 PHY_8957 ();
 sky130_fd_sc_hd__decap_3 PHY_8958 ();
 sky130_fd_sc_hd__decap_3 PHY_8959 ();
 sky130_fd_sc_hd__decap_3 PHY_8960 ();
 sky130_fd_sc_hd__decap_3 PHY_8961 ();
 sky130_fd_sc_hd__decap_3 PHY_8962 ();
 sky130_fd_sc_hd__decap_3 PHY_8963 ();
 sky130_fd_sc_hd__decap_3 PHY_8964 ();
 sky130_fd_sc_hd__decap_3 PHY_8965 ();
 sky130_fd_sc_hd__decap_3 PHY_8966 ();
 sky130_fd_sc_hd__decap_3 PHY_8967 ();
 sky130_fd_sc_hd__decap_3 PHY_8968 ();
 sky130_fd_sc_hd__decap_3 PHY_8969 ();
 sky130_fd_sc_hd__decap_3 PHY_8970 ();
 sky130_fd_sc_hd__decap_3 PHY_8971 ();
 sky130_fd_sc_hd__decap_3 PHY_8972 ();
 sky130_fd_sc_hd__decap_3 PHY_8973 ();
 sky130_fd_sc_hd__decap_3 PHY_8974 ();
 sky130_fd_sc_hd__decap_3 PHY_8975 ();
 sky130_fd_sc_hd__decap_3 PHY_8976 ();
 sky130_fd_sc_hd__decap_3 PHY_8977 ();
 sky130_fd_sc_hd__decap_3 PHY_8978 ();
 sky130_fd_sc_hd__decap_3 PHY_8979 ();
 sky130_fd_sc_hd__decap_3 PHY_8980 ();
 sky130_fd_sc_hd__decap_3 PHY_8981 ();
 sky130_fd_sc_hd__decap_3 PHY_8982 ();
 sky130_fd_sc_hd__decap_3 PHY_8983 ();
 sky130_fd_sc_hd__decap_3 PHY_8984 ();
 sky130_fd_sc_hd__decap_3 PHY_8985 ();
 sky130_fd_sc_hd__decap_3 PHY_8986 ();
 sky130_fd_sc_hd__decap_3 PHY_8987 ();
 sky130_fd_sc_hd__decap_3 PHY_8988 ();
 sky130_fd_sc_hd__decap_3 PHY_8989 ();
 sky130_fd_sc_hd__decap_3 PHY_8990 ();
 sky130_fd_sc_hd__decap_3 PHY_8991 ();
 sky130_fd_sc_hd__decap_3 PHY_8992 ();
 sky130_fd_sc_hd__decap_3 PHY_8993 ();
 sky130_fd_sc_hd__decap_3 PHY_8994 ();
 sky130_fd_sc_hd__decap_3 PHY_8995 ();
 sky130_fd_sc_hd__decap_3 PHY_8996 ();
 sky130_fd_sc_hd__decap_3 PHY_8997 ();
 sky130_fd_sc_hd__decap_3 PHY_8998 ();
 sky130_fd_sc_hd__decap_3 PHY_8999 ();
 sky130_fd_sc_hd__decap_3 PHY_9000 ();
 sky130_fd_sc_hd__decap_3 PHY_9001 ();
 sky130_fd_sc_hd__decap_3 PHY_9002 ();
 sky130_fd_sc_hd__decap_3 PHY_9003 ();
 sky130_fd_sc_hd__decap_3 PHY_9004 ();
 sky130_fd_sc_hd__decap_3 PHY_9005 ();
 sky130_fd_sc_hd__decap_3 PHY_9006 ();
 sky130_fd_sc_hd__decap_3 PHY_9007 ();
 sky130_fd_sc_hd__decap_3 PHY_9008 ();
 sky130_fd_sc_hd__decap_3 PHY_9009 ();
 sky130_fd_sc_hd__decap_3 PHY_9010 ();
 sky130_fd_sc_hd__decap_3 PHY_9011 ();
 sky130_fd_sc_hd__decap_3 PHY_9012 ();
 sky130_fd_sc_hd__decap_3 PHY_9013 ();
 sky130_fd_sc_hd__decap_3 PHY_9014 ();
 sky130_fd_sc_hd__decap_3 PHY_9015 ();
 sky130_fd_sc_hd__decap_3 PHY_9016 ();
 sky130_fd_sc_hd__decap_3 PHY_9017 ();
 sky130_fd_sc_hd__decap_3 PHY_9018 ();
 sky130_fd_sc_hd__decap_3 PHY_9019 ();
 sky130_fd_sc_hd__decap_3 PHY_9020 ();
 sky130_fd_sc_hd__decap_3 PHY_9021 ();
 sky130_fd_sc_hd__decap_3 PHY_9022 ();
 sky130_fd_sc_hd__decap_3 PHY_9023 ();
 sky130_fd_sc_hd__decap_3 PHY_9024 ();
 sky130_fd_sc_hd__decap_3 PHY_9025 ();
 sky130_fd_sc_hd__decap_3 PHY_9026 ();
 sky130_fd_sc_hd__decap_3 PHY_9027 ();
 sky130_fd_sc_hd__decap_3 PHY_9028 ();
 sky130_fd_sc_hd__decap_3 PHY_9029 ();
 sky130_fd_sc_hd__decap_3 PHY_9030 ();
 sky130_fd_sc_hd__decap_3 PHY_9031 ();
 sky130_fd_sc_hd__decap_3 PHY_9032 ();
 sky130_fd_sc_hd__decap_3 PHY_9033 ();
 sky130_fd_sc_hd__decap_3 PHY_9034 ();
 sky130_fd_sc_hd__decap_3 PHY_9035 ();
 sky130_fd_sc_hd__decap_3 PHY_9036 ();
 sky130_fd_sc_hd__decap_3 PHY_9037 ();
 sky130_fd_sc_hd__decap_3 PHY_9038 ();
 sky130_fd_sc_hd__decap_3 PHY_9039 ();
 sky130_fd_sc_hd__decap_3 PHY_9040 ();
 sky130_fd_sc_hd__decap_3 PHY_9041 ();
 sky130_fd_sc_hd__decap_3 PHY_9042 ();
 sky130_fd_sc_hd__decap_3 PHY_9043 ();
 sky130_fd_sc_hd__decap_3 PHY_9044 ();
 sky130_fd_sc_hd__decap_3 PHY_9045 ();
 sky130_fd_sc_hd__decap_3 PHY_9046 ();
 sky130_fd_sc_hd__decap_3 PHY_9047 ();
 sky130_fd_sc_hd__decap_3 PHY_9048 ();
 sky130_fd_sc_hd__decap_3 PHY_9049 ();
 sky130_fd_sc_hd__decap_3 PHY_9050 ();
 sky130_fd_sc_hd__decap_3 PHY_9051 ();
 sky130_fd_sc_hd__decap_3 PHY_9052 ();
 sky130_fd_sc_hd__decap_3 PHY_9053 ();
 sky130_fd_sc_hd__decap_3 PHY_9054 ();
 sky130_fd_sc_hd__decap_3 PHY_9055 ();
 sky130_fd_sc_hd__decap_3 PHY_9056 ();
 sky130_fd_sc_hd__decap_3 PHY_9057 ();
 sky130_fd_sc_hd__decap_3 PHY_9058 ();
 sky130_fd_sc_hd__decap_3 PHY_9059 ();
 sky130_fd_sc_hd__decap_3 PHY_9060 ();
 sky130_fd_sc_hd__decap_3 PHY_9061 ();
 sky130_fd_sc_hd__decap_3 PHY_9062 ();
 sky130_fd_sc_hd__decap_3 PHY_9063 ();
 sky130_fd_sc_hd__decap_3 PHY_9064 ();
 sky130_fd_sc_hd__decap_3 PHY_9065 ();
 sky130_fd_sc_hd__decap_3 PHY_9066 ();
 sky130_fd_sc_hd__decap_3 PHY_9067 ();
 sky130_fd_sc_hd__decap_3 PHY_9068 ();
 sky130_fd_sc_hd__decap_3 PHY_9069 ();
 sky130_fd_sc_hd__decap_3 PHY_9070 ();
 sky130_fd_sc_hd__decap_3 PHY_9071 ();
 sky130_fd_sc_hd__decap_3 PHY_9072 ();
 sky130_fd_sc_hd__decap_3 PHY_9073 ();
 sky130_fd_sc_hd__decap_3 PHY_9074 ();
 sky130_fd_sc_hd__decap_3 PHY_9075 ();
 sky130_fd_sc_hd__decap_3 PHY_9076 ();
 sky130_fd_sc_hd__decap_3 PHY_9077 ();
 sky130_fd_sc_hd__decap_3 PHY_9078 ();
 sky130_fd_sc_hd__decap_3 PHY_9079 ();
 sky130_fd_sc_hd__decap_3 PHY_9080 ();
 sky130_fd_sc_hd__decap_3 PHY_9081 ();
 sky130_fd_sc_hd__decap_3 PHY_9082 ();
 sky130_fd_sc_hd__decap_3 PHY_9083 ();
 sky130_fd_sc_hd__decap_3 PHY_9084 ();
 sky130_fd_sc_hd__decap_3 PHY_9085 ();
 sky130_fd_sc_hd__decap_3 PHY_9086 ();
 sky130_fd_sc_hd__decap_3 PHY_9087 ();
 sky130_fd_sc_hd__decap_3 PHY_9088 ();
 sky130_fd_sc_hd__decap_3 PHY_9089 ();
 sky130_fd_sc_hd__decap_3 PHY_9090 ();
 sky130_fd_sc_hd__decap_3 PHY_9091 ();
 sky130_fd_sc_hd__decap_3 PHY_9092 ();
 sky130_fd_sc_hd__decap_3 PHY_9093 ();
 sky130_fd_sc_hd__decap_3 PHY_9094 ();
 sky130_fd_sc_hd__decap_3 PHY_9095 ();
 sky130_fd_sc_hd__decap_3 PHY_9096 ();
 sky130_fd_sc_hd__decap_3 PHY_9097 ();
 sky130_fd_sc_hd__decap_3 PHY_9098 ();
 sky130_fd_sc_hd__decap_3 PHY_9099 ();
 sky130_fd_sc_hd__decap_3 PHY_9100 ();
 sky130_fd_sc_hd__decap_3 PHY_9101 ();
 sky130_fd_sc_hd__decap_3 PHY_9102 ();
 sky130_fd_sc_hd__decap_3 PHY_9103 ();
 sky130_fd_sc_hd__decap_3 PHY_9104 ();
 sky130_fd_sc_hd__decap_3 PHY_9105 ();
 sky130_fd_sc_hd__decap_3 PHY_9106 ();
 sky130_fd_sc_hd__decap_3 PHY_9107 ();
 sky130_fd_sc_hd__decap_3 PHY_9108 ();
 sky130_fd_sc_hd__decap_3 PHY_9109 ();
 sky130_fd_sc_hd__decap_3 PHY_9110 ();
 sky130_fd_sc_hd__decap_3 PHY_9111 ();
 sky130_fd_sc_hd__decap_3 PHY_9112 ();
 sky130_fd_sc_hd__decap_3 PHY_9113 ();
 sky130_fd_sc_hd__decap_3 PHY_9114 ();
 sky130_fd_sc_hd__decap_3 PHY_9115 ();
 sky130_fd_sc_hd__decap_3 PHY_9116 ();
 sky130_fd_sc_hd__decap_3 PHY_9117 ();
 sky130_fd_sc_hd__decap_3 PHY_9118 ();
 sky130_fd_sc_hd__decap_3 PHY_9119 ();
 sky130_fd_sc_hd__decap_3 PHY_9120 ();
 sky130_fd_sc_hd__decap_3 PHY_9121 ();
 sky130_fd_sc_hd__decap_3 PHY_9122 ();
 sky130_fd_sc_hd__decap_3 PHY_9123 ();
 sky130_fd_sc_hd__decap_3 PHY_9124 ();
 sky130_fd_sc_hd__decap_3 PHY_9125 ();
 sky130_fd_sc_hd__decap_3 PHY_9126 ();
 sky130_fd_sc_hd__decap_3 PHY_9127 ();
 sky130_fd_sc_hd__decap_3 PHY_9128 ();
 sky130_fd_sc_hd__decap_3 PHY_9129 ();
 sky130_fd_sc_hd__decap_3 PHY_9130 ();
 sky130_fd_sc_hd__decap_3 PHY_9131 ();
 sky130_fd_sc_hd__decap_3 PHY_9132 ();
 sky130_fd_sc_hd__decap_3 PHY_9133 ();
 sky130_fd_sc_hd__decap_3 PHY_9134 ();
 sky130_fd_sc_hd__decap_3 PHY_9135 ();
 sky130_fd_sc_hd__decap_3 PHY_9136 ();
 sky130_fd_sc_hd__decap_3 PHY_9137 ();
 sky130_fd_sc_hd__decap_3 PHY_9138 ();
 sky130_fd_sc_hd__decap_3 PHY_9139 ();
 sky130_fd_sc_hd__decap_3 PHY_9140 ();
 sky130_fd_sc_hd__decap_3 PHY_9141 ();
 sky130_fd_sc_hd__decap_3 PHY_9142 ();
 sky130_fd_sc_hd__decap_3 PHY_9143 ();
 sky130_fd_sc_hd__decap_3 PHY_9144 ();
 sky130_fd_sc_hd__decap_3 PHY_9145 ();
 sky130_fd_sc_hd__decap_3 PHY_9146 ();
 sky130_fd_sc_hd__decap_3 PHY_9147 ();
 sky130_fd_sc_hd__decap_3 PHY_9148 ();
 sky130_fd_sc_hd__decap_3 PHY_9149 ();
 sky130_fd_sc_hd__decap_3 PHY_9150 ();
 sky130_fd_sc_hd__decap_3 PHY_9151 ();
 sky130_fd_sc_hd__decap_3 PHY_9152 ();
 sky130_fd_sc_hd__decap_3 PHY_9153 ();
 sky130_fd_sc_hd__decap_3 PHY_9154 ();
 sky130_fd_sc_hd__decap_3 PHY_9155 ();
 sky130_fd_sc_hd__decap_3 PHY_9156 ();
 sky130_fd_sc_hd__decap_3 PHY_9157 ();
 sky130_fd_sc_hd__decap_3 PHY_9158 ();
 sky130_fd_sc_hd__decap_3 PHY_9159 ();
 sky130_fd_sc_hd__decap_3 PHY_9160 ();
 sky130_fd_sc_hd__decap_3 PHY_9161 ();
 sky130_fd_sc_hd__decap_3 PHY_9162 ();
 sky130_fd_sc_hd__decap_3 PHY_9163 ();
 sky130_fd_sc_hd__decap_3 PHY_9164 ();
 sky130_fd_sc_hd__decap_3 PHY_9165 ();
 sky130_fd_sc_hd__decap_3 PHY_9166 ();
 sky130_fd_sc_hd__decap_3 PHY_9167 ();
 sky130_fd_sc_hd__decap_3 PHY_9168 ();
 sky130_fd_sc_hd__decap_3 PHY_9169 ();
 sky130_fd_sc_hd__decap_3 PHY_9170 ();
 sky130_fd_sc_hd__decap_3 PHY_9171 ();
 sky130_fd_sc_hd__decap_3 PHY_9172 ();
 sky130_fd_sc_hd__decap_3 PHY_9173 ();
 sky130_fd_sc_hd__decap_3 PHY_9174 ();
 sky130_fd_sc_hd__decap_3 PHY_9175 ();
 sky130_fd_sc_hd__decap_3 PHY_9176 ();
 sky130_fd_sc_hd__decap_3 PHY_9177 ();
 sky130_fd_sc_hd__decap_3 PHY_9178 ();
 sky130_fd_sc_hd__decap_3 PHY_9179 ();
 sky130_fd_sc_hd__decap_3 PHY_9180 ();
 sky130_fd_sc_hd__decap_3 PHY_9181 ();
 sky130_fd_sc_hd__decap_3 PHY_9182 ();
 sky130_fd_sc_hd__decap_3 PHY_9183 ();
 sky130_fd_sc_hd__decap_3 PHY_9184 ();
 sky130_fd_sc_hd__decap_3 PHY_9185 ();
 sky130_fd_sc_hd__decap_3 PHY_9186 ();
 sky130_fd_sc_hd__decap_3 PHY_9187 ();
 sky130_fd_sc_hd__decap_3 PHY_9188 ();
 sky130_fd_sc_hd__decap_3 PHY_9189 ();
 sky130_fd_sc_hd__decap_3 PHY_9190 ();
 sky130_fd_sc_hd__decap_3 PHY_9191 ();
 sky130_fd_sc_hd__decap_3 PHY_9192 ();
 sky130_fd_sc_hd__decap_3 PHY_9193 ();
 sky130_fd_sc_hd__decap_3 PHY_9194 ();
 sky130_fd_sc_hd__decap_3 PHY_9195 ();
 sky130_fd_sc_hd__decap_3 PHY_9196 ();
 sky130_fd_sc_hd__decap_3 PHY_9197 ();
 sky130_fd_sc_hd__decap_3 PHY_9198 ();
 sky130_fd_sc_hd__decap_3 PHY_9199 ();
 sky130_fd_sc_hd__decap_3 PHY_9200 ();
 sky130_fd_sc_hd__decap_3 PHY_9201 ();
 sky130_fd_sc_hd__decap_3 PHY_9202 ();
 sky130_fd_sc_hd__decap_3 PHY_9203 ();
 sky130_fd_sc_hd__decap_3 PHY_9204 ();
 sky130_fd_sc_hd__decap_3 PHY_9205 ();
 sky130_fd_sc_hd__decap_3 PHY_9206 ();
 sky130_fd_sc_hd__decap_3 PHY_9207 ();
 sky130_fd_sc_hd__decap_3 PHY_9208 ();
 sky130_fd_sc_hd__decap_3 PHY_9209 ();
 sky130_fd_sc_hd__decap_3 PHY_9210 ();
 sky130_fd_sc_hd__decap_3 PHY_9211 ();
 sky130_fd_sc_hd__decap_3 PHY_9212 ();
 sky130_fd_sc_hd__decap_3 PHY_9213 ();
 sky130_fd_sc_hd__decap_3 PHY_9214 ();
 sky130_fd_sc_hd__decap_3 PHY_9215 ();
 sky130_fd_sc_hd__decap_3 PHY_9216 ();
 sky130_fd_sc_hd__decap_3 PHY_9217 ();
 sky130_fd_sc_hd__decap_3 PHY_9218 ();
 sky130_fd_sc_hd__decap_3 PHY_9219 ();
 sky130_fd_sc_hd__decap_3 PHY_9220 ();
 sky130_fd_sc_hd__decap_3 PHY_9221 ();
 sky130_fd_sc_hd__decap_3 PHY_9222 ();
 sky130_fd_sc_hd__decap_3 PHY_9223 ();
 sky130_fd_sc_hd__decap_3 PHY_9224 ();
 sky130_fd_sc_hd__decap_3 PHY_9225 ();
 sky130_fd_sc_hd__decap_3 PHY_9226 ();
 sky130_fd_sc_hd__decap_3 PHY_9227 ();
 sky130_fd_sc_hd__decap_3 PHY_9228 ();
 sky130_fd_sc_hd__decap_3 PHY_9229 ();
 sky130_fd_sc_hd__decap_3 PHY_9230 ();
 sky130_fd_sc_hd__decap_3 PHY_9231 ();
 sky130_fd_sc_hd__decap_3 PHY_9232 ();
 sky130_fd_sc_hd__decap_3 PHY_9233 ();
 sky130_fd_sc_hd__decap_3 PHY_9234 ();
 sky130_fd_sc_hd__decap_3 PHY_9235 ();
 sky130_fd_sc_hd__decap_3 PHY_9236 ();
 sky130_fd_sc_hd__decap_3 PHY_9237 ();
 sky130_fd_sc_hd__decap_3 PHY_9238 ();
 sky130_fd_sc_hd__decap_3 PHY_9239 ();
 sky130_fd_sc_hd__decap_3 PHY_9240 ();
 sky130_fd_sc_hd__decap_3 PHY_9241 ();
 sky130_fd_sc_hd__decap_3 PHY_9242 ();
 sky130_fd_sc_hd__decap_3 PHY_9243 ();
 sky130_fd_sc_hd__decap_3 PHY_9244 ();
 sky130_fd_sc_hd__decap_3 PHY_9245 ();
 sky130_fd_sc_hd__decap_3 PHY_9246 ();
 sky130_fd_sc_hd__decap_3 PHY_9247 ();
 sky130_fd_sc_hd__decap_3 PHY_9248 ();
 sky130_fd_sc_hd__decap_3 PHY_9249 ();
 sky130_fd_sc_hd__decap_3 PHY_9250 ();
 sky130_fd_sc_hd__decap_3 PHY_9251 ();
 sky130_fd_sc_hd__decap_3 PHY_9252 ();
 sky130_fd_sc_hd__decap_3 PHY_9253 ();
 sky130_fd_sc_hd__decap_3 PHY_9254 ();
 sky130_fd_sc_hd__decap_3 PHY_9255 ();
 sky130_fd_sc_hd__decap_3 PHY_9256 ();
 sky130_fd_sc_hd__decap_3 PHY_9257 ();
 sky130_fd_sc_hd__decap_3 PHY_9258 ();
 sky130_fd_sc_hd__decap_3 PHY_9259 ();
 sky130_fd_sc_hd__decap_3 PHY_9260 ();
 sky130_fd_sc_hd__decap_3 PHY_9261 ();
 sky130_fd_sc_hd__decap_3 PHY_9262 ();
 sky130_fd_sc_hd__decap_3 PHY_9263 ();
 sky130_fd_sc_hd__decap_3 PHY_9264 ();
 sky130_fd_sc_hd__decap_3 PHY_9265 ();
 sky130_fd_sc_hd__decap_3 PHY_9266 ();
 sky130_fd_sc_hd__decap_3 PHY_9267 ();
 sky130_fd_sc_hd__decap_3 PHY_9268 ();
 sky130_fd_sc_hd__decap_3 PHY_9269 ();
 sky130_fd_sc_hd__decap_3 PHY_9270 ();
 sky130_fd_sc_hd__decap_3 PHY_9271 ();
 sky130_fd_sc_hd__decap_3 PHY_9272 ();
 sky130_fd_sc_hd__decap_3 PHY_9273 ();
 sky130_fd_sc_hd__decap_3 PHY_9274 ();
 sky130_fd_sc_hd__decap_3 PHY_9275 ();
 sky130_fd_sc_hd__decap_3 PHY_9276 ();
 sky130_fd_sc_hd__decap_3 PHY_9277 ();
 sky130_fd_sc_hd__decap_3 PHY_9278 ();
 sky130_fd_sc_hd__decap_3 PHY_9279 ();
 sky130_fd_sc_hd__decap_3 PHY_9280 ();
 sky130_fd_sc_hd__decap_3 PHY_9281 ();
 sky130_fd_sc_hd__decap_3 PHY_9282 ();
 sky130_fd_sc_hd__decap_3 PHY_9283 ();
 sky130_fd_sc_hd__decap_3 PHY_9284 ();
 sky130_fd_sc_hd__decap_3 PHY_9285 ();
 sky130_fd_sc_hd__decap_3 PHY_9286 ();
 sky130_fd_sc_hd__decap_3 PHY_9287 ();
 sky130_fd_sc_hd__decap_3 PHY_9288 ();
 sky130_fd_sc_hd__decap_3 PHY_9289 ();
 sky130_fd_sc_hd__decap_3 PHY_9290 ();
 sky130_fd_sc_hd__decap_3 PHY_9291 ();
 sky130_fd_sc_hd__decap_3 PHY_9292 ();
 sky130_fd_sc_hd__decap_3 PHY_9293 ();
 sky130_fd_sc_hd__decap_3 PHY_9294 ();
 sky130_fd_sc_hd__decap_3 PHY_9295 ();
 sky130_fd_sc_hd__decap_3 PHY_9296 ();
 sky130_fd_sc_hd__decap_3 PHY_9297 ();
 sky130_fd_sc_hd__decap_3 PHY_9298 ();
 sky130_fd_sc_hd__decap_3 PHY_9299 ();
 sky130_fd_sc_hd__decap_3 PHY_9300 ();
 sky130_fd_sc_hd__decap_3 PHY_9301 ();
 sky130_fd_sc_hd__decap_3 PHY_9302 ();
 sky130_fd_sc_hd__decap_3 PHY_9303 ();
 sky130_fd_sc_hd__decap_3 PHY_9304 ();
 sky130_fd_sc_hd__decap_3 PHY_9305 ();
 sky130_fd_sc_hd__decap_3 PHY_9306 ();
 sky130_fd_sc_hd__decap_3 PHY_9307 ();
 sky130_fd_sc_hd__decap_3 PHY_9308 ();
 sky130_fd_sc_hd__decap_3 PHY_9309 ();
 sky130_fd_sc_hd__decap_3 PHY_9310 ();
 sky130_fd_sc_hd__decap_3 PHY_9311 ();
 sky130_fd_sc_hd__decap_3 PHY_9312 ();
 sky130_fd_sc_hd__decap_3 PHY_9313 ();
 sky130_fd_sc_hd__decap_3 PHY_9314 ();
 sky130_fd_sc_hd__decap_3 PHY_9315 ();
 sky130_fd_sc_hd__decap_3 PHY_9316 ();
 sky130_fd_sc_hd__decap_3 PHY_9317 ();
 sky130_fd_sc_hd__decap_3 PHY_9318 ();
 sky130_fd_sc_hd__decap_3 PHY_9319 ();
 sky130_fd_sc_hd__decap_3 PHY_9320 ();
 sky130_fd_sc_hd__decap_3 PHY_9321 ();
 sky130_fd_sc_hd__decap_3 PHY_9322 ();
 sky130_fd_sc_hd__decap_3 PHY_9323 ();
 sky130_fd_sc_hd__decap_3 PHY_9324 ();
 sky130_fd_sc_hd__decap_3 PHY_9325 ();
 sky130_fd_sc_hd__decap_3 PHY_9326 ();
 sky130_fd_sc_hd__decap_3 PHY_9327 ();
 sky130_fd_sc_hd__decap_3 PHY_9328 ();
 sky130_fd_sc_hd__decap_3 PHY_9329 ();
 sky130_fd_sc_hd__decap_3 PHY_9330 ();
 sky130_fd_sc_hd__decap_3 PHY_9331 ();
 sky130_fd_sc_hd__decap_3 PHY_9332 ();
 sky130_fd_sc_hd__decap_3 PHY_9333 ();
 sky130_fd_sc_hd__decap_3 PHY_9334 ();
 sky130_fd_sc_hd__decap_3 PHY_9335 ();
 sky130_fd_sc_hd__decap_3 PHY_9336 ();
 sky130_fd_sc_hd__decap_3 PHY_9337 ();
 sky130_fd_sc_hd__decap_3 PHY_9338 ();
 sky130_fd_sc_hd__decap_3 PHY_9339 ();
 sky130_fd_sc_hd__decap_3 PHY_9340 ();
 sky130_fd_sc_hd__decap_3 PHY_9341 ();
 sky130_fd_sc_hd__decap_3 PHY_9342 ();
 sky130_fd_sc_hd__decap_3 PHY_9343 ();
 sky130_fd_sc_hd__decap_3 PHY_9344 ();
 sky130_fd_sc_hd__decap_3 PHY_9345 ();
 sky130_fd_sc_hd__decap_3 PHY_9346 ();
 sky130_fd_sc_hd__decap_3 PHY_9347 ();
 sky130_fd_sc_hd__decap_3 PHY_9348 ();
 sky130_fd_sc_hd__decap_3 PHY_9349 ();
 sky130_fd_sc_hd__decap_3 PHY_9350 ();
 sky130_fd_sc_hd__decap_3 PHY_9351 ();
 sky130_fd_sc_hd__decap_3 PHY_9352 ();
 sky130_fd_sc_hd__decap_3 PHY_9353 ();
 sky130_fd_sc_hd__decap_3 PHY_9354 ();
 sky130_fd_sc_hd__decap_3 PHY_9355 ();
 sky130_fd_sc_hd__decap_3 PHY_9356 ();
 sky130_fd_sc_hd__decap_3 PHY_9357 ();
 sky130_fd_sc_hd__decap_3 PHY_9358 ();
 sky130_fd_sc_hd__decap_3 PHY_9359 ();
 sky130_fd_sc_hd__decap_3 PHY_9360 ();
 sky130_fd_sc_hd__decap_3 PHY_9361 ();
 sky130_fd_sc_hd__decap_3 PHY_9362 ();
 sky130_fd_sc_hd__decap_3 PHY_9363 ();
 sky130_fd_sc_hd__decap_3 PHY_9364 ();
 sky130_fd_sc_hd__decap_3 PHY_9365 ();
 sky130_fd_sc_hd__decap_3 PHY_9366 ();
 sky130_fd_sc_hd__decap_3 PHY_9367 ();
 sky130_fd_sc_hd__decap_3 PHY_9368 ();
 sky130_fd_sc_hd__decap_3 PHY_9369 ();
 sky130_fd_sc_hd__decap_3 PHY_9370 ();
 sky130_fd_sc_hd__decap_3 PHY_9371 ();
 sky130_fd_sc_hd__decap_3 PHY_9372 ();
 sky130_fd_sc_hd__decap_3 PHY_9373 ();
 sky130_fd_sc_hd__decap_3 PHY_9374 ();
 sky130_fd_sc_hd__decap_3 PHY_9375 ();
 sky130_fd_sc_hd__decap_3 PHY_9376 ();
 sky130_fd_sc_hd__decap_3 PHY_9377 ();
 sky130_fd_sc_hd__decap_3 PHY_9378 ();
 sky130_fd_sc_hd__decap_3 PHY_9379 ();
 sky130_fd_sc_hd__decap_3 PHY_9380 ();
 sky130_fd_sc_hd__decap_3 PHY_9381 ();
 sky130_fd_sc_hd__decap_3 PHY_9382 ();
 sky130_fd_sc_hd__decap_3 PHY_9383 ();
 sky130_fd_sc_hd__decap_3 PHY_9384 ();
 sky130_fd_sc_hd__decap_3 PHY_9385 ();
 sky130_fd_sc_hd__decap_3 PHY_9386 ();
 sky130_fd_sc_hd__decap_3 PHY_9387 ();
 sky130_fd_sc_hd__decap_3 PHY_9388 ();
 sky130_fd_sc_hd__decap_3 PHY_9389 ();
 sky130_fd_sc_hd__decap_3 PHY_9390 ();
 sky130_fd_sc_hd__decap_3 PHY_9391 ();
 sky130_fd_sc_hd__decap_3 PHY_9392 ();
 sky130_fd_sc_hd__decap_3 PHY_9393 ();
 sky130_fd_sc_hd__decap_3 PHY_9394 ();
 sky130_fd_sc_hd__decap_3 PHY_9395 ();
 sky130_fd_sc_hd__decap_3 PHY_9396 ();
 sky130_fd_sc_hd__decap_3 PHY_9397 ();
 sky130_fd_sc_hd__decap_3 PHY_9398 ();
 sky130_fd_sc_hd__decap_3 PHY_9399 ();
 sky130_fd_sc_hd__decap_3 PHY_9400 ();
 sky130_fd_sc_hd__decap_3 PHY_9401 ();
 sky130_fd_sc_hd__decap_3 PHY_9402 ();
 sky130_fd_sc_hd__decap_3 PHY_9403 ();
 sky130_fd_sc_hd__decap_3 PHY_9404 ();
 sky130_fd_sc_hd__decap_3 PHY_9405 ();
 sky130_fd_sc_hd__decap_3 PHY_9406 ();
 sky130_fd_sc_hd__decap_3 PHY_9407 ();
 sky130_fd_sc_hd__decap_3 PHY_9408 ();
 sky130_fd_sc_hd__decap_3 PHY_9409 ();
 sky130_fd_sc_hd__decap_3 PHY_9410 ();
 sky130_fd_sc_hd__decap_3 PHY_9411 ();
 sky130_fd_sc_hd__decap_3 PHY_9412 ();
 sky130_fd_sc_hd__decap_3 PHY_9413 ();
 sky130_fd_sc_hd__decap_3 PHY_9414 ();
 sky130_fd_sc_hd__decap_3 PHY_9415 ();
 sky130_fd_sc_hd__decap_3 PHY_9416 ();
 sky130_fd_sc_hd__decap_3 PHY_9417 ();
 sky130_fd_sc_hd__decap_3 PHY_9418 ();
 sky130_fd_sc_hd__decap_3 PHY_9419 ();
 sky130_fd_sc_hd__decap_3 PHY_9420 ();
 sky130_fd_sc_hd__decap_3 PHY_9421 ();
 sky130_fd_sc_hd__decap_3 PHY_9422 ();
 sky130_fd_sc_hd__decap_3 PHY_9423 ();
 sky130_fd_sc_hd__decap_3 PHY_9424 ();
 sky130_fd_sc_hd__decap_3 PHY_9425 ();
 sky130_fd_sc_hd__decap_3 PHY_9426 ();
 sky130_fd_sc_hd__decap_3 PHY_9427 ();
 sky130_fd_sc_hd__decap_3 PHY_9428 ();
 sky130_fd_sc_hd__decap_3 PHY_9429 ();
 sky130_fd_sc_hd__decap_3 PHY_9430 ();
 sky130_fd_sc_hd__decap_3 PHY_9431 ();
 sky130_fd_sc_hd__decap_3 PHY_9432 ();
 sky130_fd_sc_hd__decap_3 PHY_9433 ();
 sky130_fd_sc_hd__decap_3 PHY_9434 ();
 sky130_fd_sc_hd__decap_3 PHY_9435 ();
 sky130_fd_sc_hd__decap_3 PHY_9436 ();
 sky130_fd_sc_hd__decap_3 PHY_9437 ();
 sky130_fd_sc_hd__decap_3 PHY_9438 ();
 sky130_fd_sc_hd__decap_3 PHY_9439 ();
 sky130_fd_sc_hd__decap_3 PHY_9440 ();
 sky130_fd_sc_hd__decap_3 PHY_9441 ();
 sky130_fd_sc_hd__decap_3 PHY_9442 ();
 sky130_fd_sc_hd__decap_3 PHY_9443 ();
 sky130_fd_sc_hd__decap_3 PHY_9444 ();
 sky130_fd_sc_hd__decap_3 PHY_9445 ();
 sky130_fd_sc_hd__decap_3 PHY_9446 ();
 sky130_fd_sc_hd__decap_3 PHY_9447 ();
 sky130_fd_sc_hd__decap_3 PHY_9448 ();
 sky130_fd_sc_hd__decap_3 PHY_9449 ();
 sky130_fd_sc_hd__decap_3 PHY_9450 ();
 sky130_fd_sc_hd__decap_3 PHY_9451 ();
 sky130_fd_sc_hd__decap_3 PHY_9452 ();
 sky130_fd_sc_hd__decap_3 PHY_9453 ();
 sky130_fd_sc_hd__decap_3 PHY_9454 ();
 sky130_fd_sc_hd__decap_3 PHY_9455 ();
 sky130_fd_sc_hd__decap_3 PHY_9456 ();
 sky130_fd_sc_hd__decap_3 PHY_9457 ();
 sky130_fd_sc_hd__decap_3 PHY_9458 ();
 sky130_fd_sc_hd__decap_3 PHY_9459 ();
 sky130_fd_sc_hd__decap_3 PHY_9460 ();
 sky130_fd_sc_hd__decap_3 PHY_9461 ();
 sky130_fd_sc_hd__decap_3 PHY_9462 ();
 sky130_fd_sc_hd__decap_3 PHY_9463 ();
 sky130_fd_sc_hd__decap_3 PHY_9464 ();
 sky130_fd_sc_hd__decap_3 PHY_9465 ();
 sky130_fd_sc_hd__decap_3 PHY_9466 ();
 sky130_fd_sc_hd__decap_3 PHY_9467 ();
 sky130_fd_sc_hd__decap_3 PHY_9468 ();
 sky130_fd_sc_hd__decap_3 PHY_9469 ();
 sky130_fd_sc_hd__decap_3 PHY_9470 ();
 sky130_fd_sc_hd__decap_3 PHY_9471 ();
 sky130_fd_sc_hd__decap_3 PHY_9472 ();
 sky130_fd_sc_hd__decap_3 PHY_9473 ();
 sky130_fd_sc_hd__decap_3 PHY_9474 ();
 sky130_fd_sc_hd__decap_3 PHY_9475 ();
 sky130_fd_sc_hd__decap_3 PHY_9476 ();
 sky130_fd_sc_hd__decap_3 PHY_9477 ();
 sky130_fd_sc_hd__decap_3 PHY_9478 ();
 sky130_fd_sc_hd__decap_3 PHY_9479 ();
 sky130_fd_sc_hd__decap_3 PHY_9480 ();
 sky130_fd_sc_hd__decap_3 PHY_9481 ();
 sky130_fd_sc_hd__decap_3 PHY_9482 ();
 sky130_fd_sc_hd__decap_3 PHY_9483 ();
 sky130_fd_sc_hd__decap_3 PHY_9484 ();
 sky130_fd_sc_hd__decap_3 PHY_9485 ();
 sky130_fd_sc_hd__decap_3 PHY_9486 ();
 sky130_fd_sc_hd__decap_3 PHY_9487 ();
 sky130_fd_sc_hd__decap_3 PHY_9488 ();
 sky130_fd_sc_hd__decap_3 PHY_9489 ();
 sky130_fd_sc_hd__decap_3 PHY_9490 ();
 sky130_fd_sc_hd__decap_3 PHY_9491 ();
 sky130_fd_sc_hd__decap_3 PHY_9492 ();
 sky130_fd_sc_hd__decap_3 PHY_9493 ();
 sky130_fd_sc_hd__decap_3 PHY_9494 ();
 sky130_fd_sc_hd__decap_3 PHY_9495 ();
 sky130_fd_sc_hd__decap_3 PHY_9496 ();
 sky130_fd_sc_hd__decap_3 PHY_9497 ();
 sky130_fd_sc_hd__decap_3 PHY_9498 ();
 sky130_fd_sc_hd__decap_3 PHY_9499 ();
 sky130_fd_sc_hd__decap_3 PHY_9500 ();
 sky130_fd_sc_hd__decap_3 PHY_9501 ();
 sky130_fd_sc_hd__decap_3 PHY_9502 ();
 sky130_fd_sc_hd__decap_3 PHY_9503 ();
 sky130_fd_sc_hd__decap_3 PHY_9504 ();
 sky130_fd_sc_hd__decap_3 PHY_9505 ();
 sky130_fd_sc_hd__decap_3 PHY_9506 ();
 sky130_fd_sc_hd__decap_3 PHY_9507 ();
 sky130_fd_sc_hd__decap_3 PHY_9508 ();
 sky130_fd_sc_hd__decap_3 PHY_9509 ();
 sky130_fd_sc_hd__decap_3 PHY_9510 ();
 sky130_fd_sc_hd__decap_3 PHY_9511 ();
 sky130_fd_sc_hd__decap_3 PHY_9512 ();
 sky130_fd_sc_hd__decap_3 PHY_9513 ();
 sky130_fd_sc_hd__decap_3 PHY_9514 ();
 sky130_fd_sc_hd__decap_3 PHY_9515 ();
 sky130_fd_sc_hd__decap_3 PHY_9516 ();
 sky130_fd_sc_hd__decap_3 PHY_9517 ();
 sky130_fd_sc_hd__decap_3 PHY_9518 ();
 sky130_fd_sc_hd__decap_3 PHY_9519 ();
 sky130_fd_sc_hd__decap_3 PHY_9520 ();
 sky130_fd_sc_hd__decap_3 PHY_9521 ();
 sky130_fd_sc_hd__decap_3 PHY_9522 ();
 sky130_fd_sc_hd__decap_3 PHY_9523 ();
 sky130_fd_sc_hd__decap_3 PHY_9524 ();
 sky130_fd_sc_hd__decap_3 PHY_9525 ();
 sky130_fd_sc_hd__decap_3 PHY_9526 ();
 sky130_fd_sc_hd__decap_3 PHY_9527 ();
 sky130_fd_sc_hd__decap_3 PHY_9528 ();
 sky130_fd_sc_hd__decap_3 PHY_9529 ();
 sky130_fd_sc_hd__decap_3 PHY_9530 ();
 sky130_fd_sc_hd__decap_3 PHY_9531 ();
 sky130_fd_sc_hd__decap_3 PHY_9532 ();
 sky130_fd_sc_hd__decap_3 PHY_9533 ();
 sky130_fd_sc_hd__decap_3 PHY_9534 ();
 sky130_fd_sc_hd__decap_3 PHY_9535 ();
 sky130_fd_sc_hd__decap_3 PHY_9536 ();
 sky130_fd_sc_hd__decap_3 PHY_9537 ();
 sky130_fd_sc_hd__decap_3 PHY_9538 ();
 sky130_fd_sc_hd__decap_3 PHY_9539 ();
 sky130_fd_sc_hd__decap_3 PHY_9540 ();
 sky130_fd_sc_hd__decap_3 PHY_9541 ();
 sky130_fd_sc_hd__decap_3 PHY_9542 ();
 sky130_fd_sc_hd__decap_3 PHY_9543 ();
 sky130_fd_sc_hd__decap_3 PHY_9544 ();
 sky130_fd_sc_hd__decap_3 PHY_9545 ();
 sky130_fd_sc_hd__decap_3 PHY_9546 ();
 sky130_fd_sc_hd__decap_3 PHY_9547 ();
 sky130_fd_sc_hd__decap_3 PHY_9548 ();
 sky130_fd_sc_hd__decap_3 PHY_9549 ();
 sky130_fd_sc_hd__decap_3 PHY_9550 ();
 sky130_fd_sc_hd__decap_3 PHY_9551 ();
 sky130_fd_sc_hd__decap_3 PHY_9552 ();
 sky130_fd_sc_hd__decap_3 PHY_9553 ();
 sky130_fd_sc_hd__decap_3 PHY_9554 ();
 sky130_fd_sc_hd__decap_3 PHY_9555 ();
 sky130_fd_sc_hd__decap_3 PHY_9556 ();
 sky130_fd_sc_hd__decap_3 PHY_9557 ();
 sky130_fd_sc_hd__decap_3 PHY_9558 ();
 sky130_fd_sc_hd__decap_3 PHY_9559 ();
 sky130_fd_sc_hd__decap_3 PHY_9560 ();
 sky130_fd_sc_hd__decap_3 PHY_9561 ();
 sky130_fd_sc_hd__decap_3 PHY_9562 ();
 sky130_fd_sc_hd__decap_3 PHY_9563 ();
 sky130_fd_sc_hd__decap_3 PHY_9564 ();
 sky130_fd_sc_hd__decap_3 PHY_9565 ();
 sky130_fd_sc_hd__decap_3 PHY_9566 ();
 sky130_fd_sc_hd__decap_3 PHY_9567 ();
 sky130_fd_sc_hd__decap_3 PHY_9568 ();
 sky130_fd_sc_hd__decap_3 PHY_9569 ();
 sky130_fd_sc_hd__decap_3 PHY_9570 ();
 sky130_fd_sc_hd__decap_3 PHY_9571 ();
 sky130_fd_sc_hd__decap_3 PHY_9572 ();
 sky130_fd_sc_hd__decap_3 PHY_9573 ();
 sky130_fd_sc_hd__decap_3 PHY_9574 ();
 sky130_fd_sc_hd__decap_3 PHY_9575 ();
 sky130_fd_sc_hd__decap_3 PHY_9576 ();
 sky130_fd_sc_hd__decap_3 PHY_9577 ();
 sky130_fd_sc_hd__decap_3 PHY_9578 ();
 sky130_fd_sc_hd__decap_3 PHY_9579 ();
 sky130_fd_sc_hd__decap_3 PHY_9580 ();
 sky130_fd_sc_hd__decap_3 PHY_9581 ();
 sky130_fd_sc_hd__decap_3 PHY_9582 ();
 sky130_fd_sc_hd__decap_3 PHY_9583 ();
 sky130_fd_sc_hd__decap_3 PHY_9584 ();
 sky130_fd_sc_hd__decap_3 PHY_9585 ();
 sky130_fd_sc_hd__decap_3 PHY_9586 ();
 sky130_fd_sc_hd__decap_3 PHY_9587 ();
 sky130_fd_sc_hd__decap_3 PHY_9588 ();
 sky130_fd_sc_hd__decap_3 PHY_9589 ();
 sky130_fd_sc_hd__decap_3 PHY_9590 ();
 sky130_fd_sc_hd__decap_3 PHY_9591 ();
 sky130_fd_sc_hd__decap_3 PHY_9592 ();
 sky130_fd_sc_hd__decap_3 PHY_9593 ();
 sky130_fd_sc_hd__decap_3 PHY_9594 ();
 sky130_fd_sc_hd__decap_3 PHY_9595 ();
 sky130_fd_sc_hd__decap_3 PHY_9596 ();
 sky130_fd_sc_hd__decap_3 PHY_9597 ();
 sky130_fd_sc_hd__decap_3 PHY_9598 ();
 sky130_fd_sc_hd__decap_3 PHY_9599 ();
 sky130_fd_sc_hd__decap_3 PHY_9600 ();
 sky130_fd_sc_hd__decap_3 PHY_9601 ();
 sky130_fd_sc_hd__decap_3 PHY_9602 ();
 sky130_fd_sc_hd__decap_3 PHY_9603 ();
 sky130_fd_sc_hd__decap_3 PHY_9604 ();
 sky130_fd_sc_hd__decap_3 PHY_9605 ();
 sky130_fd_sc_hd__decap_3 PHY_9606 ();
 sky130_fd_sc_hd__decap_3 PHY_9607 ();
 sky130_fd_sc_hd__decap_3 PHY_9608 ();
 sky130_fd_sc_hd__decap_3 PHY_9609 ();
 sky130_fd_sc_hd__decap_3 PHY_9610 ();
 sky130_fd_sc_hd__decap_3 PHY_9611 ();
 sky130_fd_sc_hd__decap_3 PHY_9612 ();
 sky130_fd_sc_hd__decap_3 PHY_9613 ();
 sky130_fd_sc_hd__decap_3 PHY_9614 ();
 sky130_fd_sc_hd__decap_3 PHY_9615 ();
 sky130_fd_sc_hd__decap_3 PHY_9616 ();
 sky130_fd_sc_hd__decap_3 PHY_9617 ();
 sky130_fd_sc_hd__decap_3 PHY_9618 ();
 sky130_fd_sc_hd__decap_3 PHY_9619 ();
 sky130_fd_sc_hd__decap_3 PHY_9620 ();
 sky130_fd_sc_hd__decap_3 PHY_9621 ();
 sky130_fd_sc_hd__decap_3 PHY_9622 ();
 sky130_fd_sc_hd__decap_3 PHY_9623 ();
 sky130_fd_sc_hd__decap_3 PHY_9624 ();
 sky130_fd_sc_hd__decap_3 PHY_9625 ();
 sky130_fd_sc_hd__decap_3 PHY_9626 ();
 sky130_fd_sc_hd__decap_3 PHY_9627 ();
 sky130_fd_sc_hd__decap_3 PHY_9628 ();
 sky130_fd_sc_hd__decap_3 PHY_9629 ();
 sky130_fd_sc_hd__decap_3 PHY_9630 ();
 sky130_fd_sc_hd__decap_3 PHY_9631 ();
 sky130_fd_sc_hd__decap_3 PHY_9632 ();
 sky130_fd_sc_hd__decap_3 PHY_9633 ();
 sky130_fd_sc_hd__decap_3 PHY_9634 ();
 sky130_fd_sc_hd__decap_3 PHY_9635 ();
 sky130_fd_sc_hd__decap_3 PHY_9636 ();
 sky130_fd_sc_hd__decap_3 PHY_9637 ();
 sky130_fd_sc_hd__decap_3 PHY_9638 ();
 sky130_fd_sc_hd__decap_3 PHY_9639 ();
 sky130_fd_sc_hd__decap_3 PHY_9640 ();
 sky130_fd_sc_hd__decap_3 PHY_9641 ();
 sky130_fd_sc_hd__decap_3 PHY_9642 ();
 sky130_fd_sc_hd__decap_3 PHY_9643 ();
 sky130_fd_sc_hd__decap_3 PHY_9644 ();
 sky130_fd_sc_hd__decap_3 PHY_9645 ();
 sky130_fd_sc_hd__decap_3 PHY_9646 ();
 sky130_fd_sc_hd__decap_3 PHY_9647 ();
 sky130_fd_sc_hd__decap_3 PHY_9648 ();
 sky130_fd_sc_hd__decap_3 PHY_9649 ();
 sky130_fd_sc_hd__decap_3 PHY_9650 ();
 sky130_fd_sc_hd__decap_3 PHY_9651 ();
 sky130_fd_sc_hd__decap_3 PHY_9652 ();
 sky130_fd_sc_hd__decap_3 PHY_9653 ();
 sky130_fd_sc_hd__decap_3 PHY_9654 ();
 sky130_fd_sc_hd__decap_3 PHY_9655 ();
 sky130_fd_sc_hd__decap_3 PHY_9656 ();
 sky130_fd_sc_hd__decap_3 PHY_9657 ();
 sky130_fd_sc_hd__decap_3 PHY_9658 ();
 sky130_fd_sc_hd__decap_3 PHY_9659 ();
 sky130_fd_sc_hd__decap_3 PHY_9660 ();
 sky130_fd_sc_hd__decap_3 PHY_9661 ();
 sky130_fd_sc_hd__decap_3 PHY_9662 ();
 sky130_fd_sc_hd__decap_3 PHY_9663 ();
 sky130_fd_sc_hd__decap_3 PHY_9664 ();
 sky130_fd_sc_hd__decap_3 PHY_9665 ();
 sky130_fd_sc_hd__decap_3 PHY_9666 ();
 sky130_fd_sc_hd__decap_3 PHY_9667 ();
 sky130_fd_sc_hd__decap_3 PHY_9668 ();
 sky130_fd_sc_hd__decap_3 PHY_9669 ();
 sky130_fd_sc_hd__decap_3 PHY_9670 ();
 sky130_fd_sc_hd__decap_3 PHY_9671 ();
 sky130_fd_sc_hd__decap_3 PHY_9672 ();
 sky130_fd_sc_hd__decap_3 PHY_9673 ();
 sky130_fd_sc_hd__decap_3 PHY_9674 ();
 sky130_fd_sc_hd__decap_3 PHY_9675 ();
 sky130_fd_sc_hd__decap_3 PHY_9676 ();
 sky130_fd_sc_hd__decap_3 PHY_9677 ();
 sky130_fd_sc_hd__decap_3 PHY_9678 ();
 sky130_fd_sc_hd__decap_3 PHY_9679 ();
 sky130_fd_sc_hd__decap_3 PHY_9680 ();
 sky130_fd_sc_hd__decap_3 PHY_9681 ();
 sky130_fd_sc_hd__decap_3 PHY_9682 ();
 sky130_fd_sc_hd__decap_3 PHY_9683 ();
 sky130_fd_sc_hd__decap_3 PHY_9684 ();
 sky130_fd_sc_hd__decap_3 PHY_9685 ();
 sky130_fd_sc_hd__decap_3 PHY_9686 ();
 sky130_fd_sc_hd__decap_3 PHY_9687 ();
 sky130_fd_sc_hd__decap_3 PHY_9688 ();
 sky130_fd_sc_hd__decap_3 PHY_9689 ();
 sky130_fd_sc_hd__decap_3 PHY_9690 ();
 sky130_fd_sc_hd__decap_3 PHY_9691 ();
 sky130_fd_sc_hd__decap_3 PHY_9692 ();
 sky130_fd_sc_hd__decap_3 PHY_9693 ();
 sky130_fd_sc_hd__decap_3 PHY_9694 ();
 sky130_fd_sc_hd__decap_3 PHY_9695 ();
 sky130_fd_sc_hd__decap_3 PHY_9696 ();
 sky130_fd_sc_hd__decap_3 PHY_9697 ();
 sky130_fd_sc_hd__decap_3 PHY_9698 ();
 sky130_fd_sc_hd__decap_3 PHY_9699 ();
 sky130_fd_sc_hd__decap_3 PHY_9700 ();
 sky130_fd_sc_hd__decap_3 PHY_9701 ();
 sky130_fd_sc_hd__decap_3 PHY_9702 ();
 sky130_fd_sc_hd__decap_3 PHY_9703 ();
 sky130_fd_sc_hd__decap_3 PHY_9704 ();
 sky130_fd_sc_hd__decap_3 PHY_9705 ();
 sky130_fd_sc_hd__decap_3 PHY_9706 ();
 sky130_fd_sc_hd__decap_3 PHY_9707 ();
 sky130_fd_sc_hd__decap_3 PHY_9708 ();
 sky130_fd_sc_hd__decap_3 PHY_9709 ();
 sky130_fd_sc_hd__decap_3 PHY_9710 ();
 sky130_fd_sc_hd__decap_3 PHY_9711 ();
 sky130_fd_sc_hd__decap_3 PHY_9712 ();
 sky130_fd_sc_hd__decap_3 PHY_9713 ();
 sky130_fd_sc_hd__decap_3 PHY_9714 ();
 sky130_fd_sc_hd__decap_3 PHY_9715 ();
 sky130_fd_sc_hd__decap_3 PHY_9716 ();
 sky130_fd_sc_hd__decap_3 PHY_9717 ();
 sky130_fd_sc_hd__decap_3 PHY_9718 ();
 sky130_fd_sc_hd__decap_3 PHY_9719 ();
 sky130_fd_sc_hd__decap_3 PHY_9720 ();
 sky130_fd_sc_hd__decap_3 PHY_9721 ();
 sky130_fd_sc_hd__decap_3 PHY_9722 ();
 sky130_fd_sc_hd__decap_3 PHY_9723 ();
 sky130_fd_sc_hd__decap_3 PHY_9724 ();
 sky130_fd_sc_hd__decap_3 PHY_9725 ();
 sky130_fd_sc_hd__decap_3 PHY_9726 ();
 sky130_fd_sc_hd__decap_3 PHY_9727 ();
 sky130_fd_sc_hd__decap_3 PHY_9728 ();
 sky130_fd_sc_hd__decap_3 PHY_9729 ();
 sky130_fd_sc_hd__decap_3 PHY_9730 ();
 sky130_fd_sc_hd__decap_3 PHY_9731 ();
 sky130_fd_sc_hd__decap_3 PHY_9732 ();
 sky130_fd_sc_hd__decap_3 PHY_9733 ();
 sky130_fd_sc_hd__decap_3 PHY_9734 ();
 sky130_fd_sc_hd__decap_3 PHY_9735 ();
 sky130_fd_sc_hd__decap_3 PHY_9736 ();
 sky130_fd_sc_hd__decap_3 PHY_9737 ();
 sky130_fd_sc_hd__decap_3 PHY_9738 ();
 sky130_fd_sc_hd__decap_3 PHY_9739 ();
 sky130_fd_sc_hd__decap_3 PHY_9740 ();
 sky130_fd_sc_hd__decap_3 PHY_9741 ();
 sky130_fd_sc_hd__decap_3 PHY_9742 ();
 sky130_fd_sc_hd__decap_3 PHY_9743 ();
 sky130_fd_sc_hd__decap_3 PHY_9744 ();
 sky130_fd_sc_hd__decap_3 PHY_9745 ();
 sky130_fd_sc_hd__decap_3 PHY_9746 ();
 sky130_fd_sc_hd__decap_3 PHY_9747 ();
 sky130_fd_sc_hd__decap_3 PHY_9748 ();
 sky130_fd_sc_hd__decap_3 PHY_9749 ();
 sky130_fd_sc_hd__decap_3 PHY_9750 ();
 sky130_fd_sc_hd__decap_3 PHY_9751 ();
 sky130_fd_sc_hd__decap_3 PHY_9752 ();
 sky130_fd_sc_hd__decap_3 PHY_9753 ();
 sky130_fd_sc_hd__decap_3 PHY_9754 ();
 sky130_fd_sc_hd__decap_3 PHY_9755 ();
 sky130_fd_sc_hd__decap_3 PHY_9756 ();
 sky130_fd_sc_hd__decap_3 PHY_9757 ();
 sky130_fd_sc_hd__decap_3 PHY_9758 ();
 sky130_fd_sc_hd__decap_3 PHY_9759 ();
 sky130_fd_sc_hd__decap_3 PHY_9760 ();
 sky130_fd_sc_hd__decap_3 PHY_9761 ();
 sky130_fd_sc_hd__decap_3 PHY_9762 ();
 sky130_fd_sc_hd__decap_3 PHY_9763 ();
 sky130_fd_sc_hd__decap_3 PHY_9764 ();
 sky130_fd_sc_hd__decap_3 PHY_9765 ();
 sky130_fd_sc_hd__decap_3 PHY_9766 ();
 sky130_fd_sc_hd__decap_3 PHY_9767 ();
 sky130_fd_sc_hd__decap_3 PHY_9768 ();
 sky130_fd_sc_hd__decap_3 PHY_9769 ();
 sky130_fd_sc_hd__decap_3 PHY_9770 ();
 sky130_fd_sc_hd__decap_3 PHY_9771 ();
 sky130_fd_sc_hd__decap_3 PHY_9772 ();
 sky130_fd_sc_hd__decap_3 PHY_9773 ();
 sky130_fd_sc_hd__decap_3 PHY_9774 ();
 sky130_fd_sc_hd__decap_3 PHY_9775 ();
 sky130_fd_sc_hd__decap_3 PHY_9776 ();
 sky130_fd_sc_hd__decap_3 PHY_9777 ();
 sky130_fd_sc_hd__decap_3 PHY_9778 ();
 sky130_fd_sc_hd__decap_3 PHY_9779 ();
 sky130_fd_sc_hd__decap_3 PHY_9780 ();
 sky130_fd_sc_hd__decap_3 PHY_9781 ();
 sky130_fd_sc_hd__decap_3 PHY_9782 ();
 sky130_fd_sc_hd__decap_3 PHY_9783 ();
 sky130_fd_sc_hd__decap_3 PHY_9784 ();
 sky130_fd_sc_hd__decap_3 PHY_9785 ();
 sky130_fd_sc_hd__decap_3 PHY_9786 ();
 sky130_fd_sc_hd__decap_3 PHY_9787 ();
 sky130_fd_sc_hd__decap_3 PHY_9788 ();
 sky130_fd_sc_hd__decap_3 PHY_9789 ();
 sky130_fd_sc_hd__decap_3 PHY_9790 ();
 sky130_fd_sc_hd__decap_3 PHY_9791 ();
 sky130_fd_sc_hd__decap_3 PHY_9792 ();
 sky130_fd_sc_hd__decap_3 PHY_9793 ();
 sky130_fd_sc_hd__decap_3 PHY_9794 ();
 sky130_fd_sc_hd__decap_3 PHY_9795 ();
 sky130_fd_sc_hd__decap_3 PHY_9796 ();
 sky130_fd_sc_hd__decap_3 PHY_9797 ();
 sky130_fd_sc_hd__decap_3 PHY_9798 ();
 sky130_fd_sc_hd__decap_3 PHY_9799 ();
 sky130_fd_sc_hd__decap_3 PHY_9800 ();
 sky130_fd_sc_hd__decap_3 PHY_9801 ();
 sky130_fd_sc_hd__decap_3 PHY_9802 ();
 sky130_fd_sc_hd__decap_3 PHY_9803 ();
 sky130_fd_sc_hd__decap_3 PHY_9804 ();
 sky130_fd_sc_hd__decap_3 PHY_9805 ();
 sky130_fd_sc_hd__decap_3 PHY_9806 ();
 sky130_fd_sc_hd__decap_3 PHY_9807 ();
 sky130_fd_sc_hd__decap_3 PHY_9808 ();
 sky130_fd_sc_hd__decap_3 PHY_9809 ();
 sky130_fd_sc_hd__decap_3 PHY_9810 ();
 sky130_fd_sc_hd__decap_3 PHY_9811 ();
 sky130_fd_sc_hd__decap_3 PHY_9812 ();
 sky130_fd_sc_hd__decap_3 PHY_9813 ();
 sky130_fd_sc_hd__decap_3 PHY_9814 ();
 sky130_fd_sc_hd__decap_3 PHY_9815 ();
 sky130_fd_sc_hd__decap_3 PHY_9816 ();
 sky130_fd_sc_hd__decap_3 PHY_9817 ();
 sky130_fd_sc_hd__decap_3 PHY_9818 ();
 sky130_fd_sc_hd__decap_3 PHY_9819 ();
 sky130_fd_sc_hd__decap_3 PHY_9820 ();
 sky130_fd_sc_hd__decap_3 PHY_9821 ();
 sky130_fd_sc_hd__decap_3 PHY_9822 ();
 sky130_fd_sc_hd__decap_3 PHY_9823 ();
 sky130_fd_sc_hd__decap_3 PHY_9824 ();
 sky130_fd_sc_hd__decap_3 PHY_9825 ();
 sky130_fd_sc_hd__decap_3 PHY_9826 ();
 sky130_fd_sc_hd__decap_3 PHY_9827 ();
 sky130_fd_sc_hd__decap_3 PHY_9828 ();
 sky130_fd_sc_hd__decap_3 PHY_9829 ();
 sky130_fd_sc_hd__decap_3 PHY_9830 ();
 sky130_fd_sc_hd__decap_3 PHY_9831 ();
 sky130_fd_sc_hd__decap_3 PHY_9832 ();
 sky130_fd_sc_hd__decap_3 PHY_9833 ();
 sky130_fd_sc_hd__decap_3 PHY_9834 ();
 sky130_fd_sc_hd__decap_3 PHY_9835 ();
 sky130_fd_sc_hd__decap_3 PHY_9836 ();
 sky130_fd_sc_hd__decap_3 PHY_9837 ();
 sky130_fd_sc_hd__decap_3 PHY_9838 ();
 sky130_fd_sc_hd__decap_3 PHY_9839 ();
 sky130_fd_sc_hd__decap_3 PHY_9840 ();
 sky130_fd_sc_hd__decap_3 PHY_9841 ();
 sky130_fd_sc_hd__decap_3 PHY_9842 ();
 sky130_fd_sc_hd__decap_3 PHY_9843 ();
 sky130_fd_sc_hd__decap_3 PHY_9844 ();
 sky130_fd_sc_hd__decap_3 PHY_9845 ();
 sky130_fd_sc_hd__decap_3 PHY_9846 ();
 sky130_fd_sc_hd__decap_3 PHY_9847 ();
 sky130_fd_sc_hd__decap_3 PHY_9848 ();
 sky130_fd_sc_hd__decap_3 PHY_9849 ();
 sky130_fd_sc_hd__decap_3 PHY_9850 ();
 sky130_fd_sc_hd__decap_3 PHY_9851 ();
 sky130_fd_sc_hd__decap_3 PHY_9852 ();
 sky130_fd_sc_hd__decap_3 PHY_9853 ();
 sky130_fd_sc_hd__decap_3 PHY_9854 ();
 sky130_fd_sc_hd__decap_3 PHY_9855 ();
 sky130_fd_sc_hd__decap_3 PHY_9856 ();
 sky130_fd_sc_hd__decap_3 PHY_9857 ();
 sky130_fd_sc_hd__decap_3 PHY_9858 ();
 sky130_fd_sc_hd__decap_3 PHY_9859 ();
 sky130_fd_sc_hd__decap_3 PHY_9860 ();
 sky130_fd_sc_hd__decap_3 PHY_9861 ();
 sky130_fd_sc_hd__decap_3 PHY_9862 ();
 sky130_fd_sc_hd__decap_3 PHY_9863 ();
 sky130_fd_sc_hd__decap_3 PHY_9864 ();
 sky130_fd_sc_hd__decap_3 PHY_9865 ();
 sky130_fd_sc_hd__decap_3 PHY_9866 ();
 sky130_fd_sc_hd__decap_3 PHY_9867 ();
 sky130_fd_sc_hd__decap_3 PHY_9868 ();
 sky130_fd_sc_hd__decap_3 PHY_9869 ();
 sky130_fd_sc_hd__decap_3 PHY_9870 ();
 sky130_fd_sc_hd__decap_3 PHY_9871 ();
 sky130_fd_sc_hd__decap_3 PHY_9872 ();
 sky130_fd_sc_hd__decap_3 PHY_9873 ();
 sky130_fd_sc_hd__decap_3 PHY_9874 ();
 sky130_fd_sc_hd__decap_3 PHY_9875 ();
 sky130_fd_sc_hd__decap_3 PHY_9876 ();
 sky130_fd_sc_hd__decap_3 PHY_9877 ();
 sky130_fd_sc_hd__decap_3 PHY_9878 ();
 sky130_fd_sc_hd__decap_3 PHY_9879 ();
 sky130_fd_sc_hd__decap_3 PHY_9880 ();
 sky130_fd_sc_hd__decap_3 PHY_9881 ();
 sky130_fd_sc_hd__decap_3 PHY_9882 ();
 sky130_fd_sc_hd__decap_3 PHY_9883 ();
 sky130_fd_sc_hd__decap_3 PHY_9884 ();
 sky130_fd_sc_hd__decap_3 PHY_9885 ();
 sky130_fd_sc_hd__decap_3 PHY_9886 ();
 sky130_fd_sc_hd__decap_3 PHY_9887 ();
 sky130_fd_sc_hd__decap_3 PHY_9888 ();
 sky130_fd_sc_hd__decap_3 PHY_9889 ();
 sky130_fd_sc_hd__decap_3 PHY_9890 ();
 sky130_fd_sc_hd__decap_3 PHY_9891 ();
 sky130_fd_sc_hd__decap_3 PHY_9892 ();
 sky130_fd_sc_hd__decap_3 PHY_9893 ();
 sky130_fd_sc_hd__decap_3 PHY_9894 ();
 sky130_fd_sc_hd__decap_3 PHY_9895 ();
 sky130_fd_sc_hd__decap_3 PHY_9896 ();
 sky130_fd_sc_hd__decap_3 PHY_9897 ();
 sky130_fd_sc_hd__decap_3 PHY_9898 ();
 sky130_fd_sc_hd__decap_3 PHY_9899 ();
 sky130_fd_sc_hd__decap_3 PHY_9900 ();
 sky130_fd_sc_hd__decap_3 PHY_9901 ();
 sky130_fd_sc_hd__decap_3 PHY_9902 ();
 sky130_fd_sc_hd__decap_3 PHY_9903 ();
 sky130_fd_sc_hd__decap_3 PHY_9904 ();
 sky130_fd_sc_hd__decap_3 PHY_9905 ();
 sky130_fd_sc_hd__decap_3 PHY_9906 ();
 sky130_fd_sc_hd__decap_3 PHY_9907 ();
 sky130_fd_sc_hd__decap_3 PHY_9908 ();
 sky130_fd_sc_hd__decap_3 PHY_9909 ();
 sky130_fd_sc_hd__decap_3 PHY_9910 ();
 sky130_fd_sc_hd__decap_3 PHY_9911 ();
 sky130_fd_sc_hd__decap_3 PHY_9912 ();
 sky130_fd_sc_hd__decap_3 PHY_9913 ();
 sky130_fd_sc_hd__decap_3 PHY_9914 ();
 sky130_fd_sc_hd__decap_3 PHY_9915 ();
 sky130_fd_sc_hd__decap_3 PHY_9916 ();
 sky130_fd_sc_hd__decap_3 PHY_9917 ();
 sky130_fd_sc_hd__decap_3 PHY_9918 ();
 sky130_fd_sc_hd__decap_3 PHY_9919 ();
 sky130_fd_sc_hd__decap_3 PHY_9920 ();
 sky130_fd_sc_hd__decap_3 PHY_9921 ();
 sky130_fd_sc_hd__decap_3 PHY_9922 ();
 sky130_fd_sc_hd__decap_3 PHY_9923 ();
 sky130_fd_sc_hd__decap_3 PHY_9924 ();
 sky130_fd_sc_hd__decap_3 PHY_9925 ();
 sky130_fd_sc_hd__decap_3 PHY_9926 ();
 sky130_fd_sc_hd__decap_3 PHY_9927 ();
 sky130_fd_sc_hd__decap_3 PHY_9928 ();
 sky130_fd_sc_hd__decap_3 PHY_9929 ();
 sky130_fd_sc_hd__decap_3 PHY_9930 ();
 sky130_fd_sc_hd__decap_3 PHY_9931 ();
 sky130_fd_sc_hd__decap_3 PHY_9932 ();
 sky130_fd_sc_hd__decap_3 PHY_9933 ();
 sky130_fd_sc_hd__decap_3 PHY_9934 ();
 sky130_fd_sc_hd__decap_3 PHY_9935 ();
 sky130_fd_sc_hd__decap_3 PHY_9936 ();
 sky130_fd_sc_hd__decap_3 PHY_9937 ();
 sky130_fd_sc_hd__decap_3 PHY_9938 ();
 sky130_fd_sc_hd__decap_3 PHY_9939 ();
 sky130_fd_sc_hd__decap_3 PHY_9940 ();
 sky130_fd_sc_hd__decap_3 PHY_9941 ();
 sky130_fd_sc_hd__decap_3 PHY_9942 ();
 sky130_fd_sc_hd__decap_3 PHY_9943 ();
 sky130_fd_sc_hd__decap_3 PHY_9944 ();
 sky130_fd_sc_hd__decap_3 PHY_9945 ();
 sky130_fd_sc_hd__decap_3 PHY_9946 ();
 sky130_fd_sc_hd__decap_3 PHY_9947 ();
 sky130_fd_sc_hd__decap_3 PHY_9948 ();
 sky130_fd_sc_hd__decap_3 PHY_9949 ();
 sky130_fd_sc_hd__decap_3 PHY_9950 ();
 sky130_fd_sc_hd__decap_3 PHY_9951 ();
 sky130_fd_sc_hd__decap_3 PHY_9952 ();
 sky130_fd_sc_hd__decap_3 PHY_9953 ();
 sky130_fd_sc_hd__decap_3 PHY_9954 ();
 sky130_fd_sc_hd__decap_3 PHY_9955 ();
 sky130_fd_sc_hd__decap_3 PHY_9956 ();
 sky130_fd_sc_hd__decap_3 PHY_9957 ();
 sky130_fd_sc_hd__decap_3 PHY_9958 ();
 sky130_fd_sc_hd__decap_3 PHY_9959 ();
 sky130_fd_sc_hd__decap_3 PHY_9960 ();
 sky130_fd_sc_hd__decap_3 PHY_9961 ();
 sky130_fd_sc_hd__decap_3 PHY_9962 ();
 sky130_fd_sc_hd__decap_3 PHY_9963 ();
 sky130_fd_sc_hd__decap_3 PHY_9964 ();
 sky130_fd_sc_hd__decap_3 PHY_9965 ();
 sky130_fd_sc_hd__decap_3 PHY_9966 ();
 sky130_fd_sc_hd__decap_3 PHY_9967 ();
 sky130_fd_sc_hd__decap_3 PHY_9968 ();
 sky130_fd_sc_hd__decap_3 PHY_9969 ();
 sky130_fd_sc_hd__decap_3 PHY_9970 ();
 sky130_fd_sc_hd__decap_3 PHY_9971 ();
 sky130_fd_sc_hd__decap_3 PHY_9972 ();
 sky130_fd_sc_hd__decap_3 PHY_9973 ();
 sky130_fd_sc_hd__decap_3 PHY_9974 ();
 sky130_fd_sc_hd__decap_3 PHY_9975 ();
 sky130_fd_sc_hd__decap_3 PHY_9976 ();
 sky130_fd_sc_hd__decap_3 PHY_9977 ();
 sky130_fd_sc_hd__decap_3 PHY_9978 ();
 sky130_fd_sc_hd__decap_3 PHY_9979 ();
 sky130_fd_sc_hd__decap_3 PHY_9980 ();
 sky130_fd_sc_hd__decap_3 PHY_9981 ();
 sky130_fd_sc_hd__decap_3 PHY_9982 ();
 sky130_fd_sc_hd__decap_3 PHY_9983 ();
 sky130_fd_sc_hd__decap_3 PHY_9984 ();
 sky130_fd_sc_hd__decap_3 PHY_9985 ();
 sky130_fd_sc_hd__decap_3 PHY_9986 ();
 sky130_fd_sc_hd__decap_3 PHY_9987 ();
 sky130_fd_sc_hd__decap_3 PHY_9988 ();
 sky130_fd_sc_hd__decap_3 PHY_9989 ();
 sky130_fd_sc_hd__decap_3 PHY_9990 ();
 sky130_fd_sc_hd__decap_3 PHY_9991 ();
 sky130_fd_sc_hd__decap_3 PHY_9992 ();
 sky130_fd_sc_hd__decap_3 PHY_9993 ();
 sky130_fd_sc_hd__decap_3 PHY_9994 ();
 sky130_fd_sc_hd__decap_3 PHY_9995 ();
 sky130_fd_sc_hd__decap_3 PHY_9996 ();
 sky130_fd_sc_hd__decap_3 PHY_9997 ();
 sky130_fd_sc_hd__decap_3 PHY_9998 ();
 sky130_fd_sc_hd__decap_3 PHY_9999 ();
 sky130_fd_sc_hd__decap_3 PHY_10000 ();
 sky130_fd_sc_hd__decap_3 PHY_10001 ();
 sky130_fd_sc_hd__decap_3 PHY_10002 ();
 sky130_fd_sc_hd__decap_3 PHY_10003 ();
 sky130_fd_sc_hd__decap_3 PHY_10004 ();
 sky130_fd_sc_hd__decap_3 PHY_10005 ();
 sky130_fd_sc_hd__decap_3 PHY_10006 ();
 sky130_fd_sc_hd__decap_3 PHY_10007 ();
 sky130_fd_sc_hd__decap_3 PHY_10008 ();
 sky130_fd_sc_hd__decap_3 PHY_10009 ();
 sky130_fd_sc_hd__decap_3 PHY_10010 ();
 sky130_fd_sc_hd__decap_3 PHY_10011 ();
 sky130_fd_sc_hd__decap_3 PHY_10012 ();
 sky130_fd_sc_hd__decap_3 PHY_10013 ();
 sky130_fd_sc_hd__decap_3 PHY_10014 ();
 sky130_fd_sc_hd__decap_3 PHY_10015 ();
 sky130_fd_sc_hd__decap_3 PHY_10016 ();
 sky130_fd_sc_hd__decap_3 PHY_10017 ();
 sky130_fd_sc_hd__decap_3 PHY_10018 ();
 sky130_fd_sc_hd__decap_3 PHY_10019 ();
 sky130_fd_sc_hd__decap_3 PHY_10020 ();
 sky130_fd_sc_hd__decap_3 PHY_10021 ();
 sky130_fd_sc_hd__decap_3 PHY_10022 ();
 sky130_fd_sc_hd__decap_3 PHY_10023 ();
 sky130_fd_sc_hd__decap_3 PHY_10024 ();
 sky130_fd_sc_hd__decap_3 PHY_10025 ();
 sky130_fd_sc_hd__decap_3 PHY_10026 ();
 sky130_fd_sc_hd__decap_3 PHY_10027 ();
 sky130_fd_sc_hd__decap_3 PHY_10028 ();
 sky130_fd_sc_hd__decap_3 PHY_10029 ();
 sky130_fd_sc_hd__decap_3 PHY_10030 ();
 sky130_fd_sc_hd__decap_3 PHY_10031 ();
 sky130_fd_sc_hd__decap_3 PHY_10032 ();
 sky130_fd_sc_hd__decap_3 PHY_10033 ();
 sky130_fd_sc_hd__decap_3 PHY_10034 ();
 sky130_fd_sc_hd__decap_3 PHY_10035 ();
 sky130_fd_sc_hd__decap_3 PHY_10036 ();
 sky130_fd_sc_hd__decap_3 PHY_10037 ();
 sky130_fd_sc_hd__decap_3 PHY_10038 ();
 sky130_fd_sc_hd__decap_3 PHY_10039 ();
 sky130_fd_sc_hd__decap_3 PHY_10040 ();
 sky130_fd_sc_hd__decap_3 PHY_10041 ();
 sky130_fd_sc_hd__decap_3 PHY_10042 ();
 sky130_fd_sc_hd__decap_3 PHY_10043 ();
 sky130_fd_sc_hd__decap_3 PHY_10044 ();
 sky130_fd_sc_hd__decap_3 PHY_10045 ();
 sky130_fd_sc_hd__decap_3 PHY_10046 ();
 sky130_fd_sc_hd__decap_3 PHY_10047 ();
 sky130_fd_sc_hd__decap_3 PHY_10048 ();
 sky130_fd_sc_hd__decap_3 PHY_10049 ();
 sky130_fd_sc_hd__decap_3 PHY_10050 ();
 sky130_fd_sc_hd__decap_3 PHY_10051 ();
 sky130_fd_sc_hd__decap_3 PHY_10052 ();
 sky130_fd_sc_hd__decap_3 PHY_10053 ();
 sky130_fd_sc_hd__decap_3 PHY_10054 ();
 sky130_fd_sc_hd__decap_3 PHY_10055 ();
 sky130_fd_sc_hd__decap_3 PHY_10056 ();
 sky130_fd_sc_hd__decap_3 PHY_10057 ();
 sky130_fd_sc_hd__decap_3 PHY_10058 ();
 sky130_fd_sc_hd__decap_3 PHY_10059 ();
 sky130_fd_sc_hd__decap_3 PHY_10060 ();
 sky130_fd_sc_hd__decap_3 PHY_10061 ();
 sky130_fd_sc_hd__decap_3 PHY_10062 ();
 sky130_fd_sc_hd__decap_3 PHY_10063 ();
 sky130_fd_sc_hd__decap_3 PHY_10064 ();
 sky130_fd_sc_hd__decap_3 PHY_10065 ();
 sky130_fd_sc_hd__decap_3 PHY_10066 ();
 sky130_fd_sc_hd__decap_3 PHY_10067 ();
 sky130_fd_sc_hd__decap_3 PHY_10068 ();
 sky130_fd_sc_hd__decap_3 PHY_10069 ();
 sky130_fd_sc_hd__decap_3 PHY_10070 ();
 sky130_fd_sc_hd__decap_3 PHY_10071 ();
 sky130_fd_sc_hd__decap_3 PHY_10072 ();
 sky130_fd_sc_hd__decap_3 PHY_10073 ();
 sky130_fd_sc_hd__decap_3 PHY_10074 ();
 sky130_fd_sc_hd__decap_3 PHY_10075 ();
 sky130_fd_sc_hd__decap_3 PHY_10076 ();
 sky130_fd_sc_hd__decap_3 PHY_10077 ();
 sky130_fd_sc_hd__decap_3 PHY_10078 ();
 sky130_fd_sc_hd__decap_3 PHY_10079 ();
 sky130_fd_sc_hd__decap_3 PHY_10080 ();
 sky130_fd_sc_hd__decap_3 PHY_10081 ();
 sky130_fd_sc_hd__decap_3 PHY_10082 ();
 sky130_fd_sc_hd__decap_3 PHY_10083 ();
 sky130_fd_sc_hd__decap_3 PHY_10084 ();
 sky130_fd_sc_hd__decap_3 PHY_10085 ();
 sky130_fd_sc_hd__decap_3 PHY_10086 ();
 sky130_fd_sc_hd__decap_3 PHY_10087 ();
 sky130_fd_sc_hd__decap_3 PHY_10088 ();
 sky130_fd_sc_hd__decap_3 PHY_10089 ();
 sky130_fd_sc_hd__decap_3 PHY_10090 ();
 sky130_fd_sc_hd__decap_3 PHY_10091 ();
 sky130_fd_sc_hd__decap_3 PHY_10092 ();
 sky130_fd_sc_hd__decap_3 PHY_10093 ();
 sky130_fd_sc_hd__decap_3 PHY_10094 ();
 sky130_fd_sc_hd__decap_3 PHY_10095 ();
 sky130_fd_sc_hd__decap_3 PHY_10096 ();
 sky130_fd_sc_hd__decap_3 PHY_10097 ();
 sky130_fd_sc_hd__decap_3 PHY_10098 ();
 sky130_fd_sc_hd__decap_3 PHY_10099 ();
 sky130_fd_sc_hd__decap_3 PHY_10100 ();
 sky130_fd_sc_hd__decap_3 PHY_10101 ();
 sky130_fd_sc_hd__decap_3 PHY_10102 ();
 sky130_fd_sc_hd__decap_3 PHY_10103 ();
 sky130_fd_sc_hd__decap_3 PHY_10104 ();
 sky130_fd_sc_hd__decap_3 PHY_10105 ();
 sky130_fd_sc_hd__decap_3 PHY_10106 ();
 sky130_fd_sc_hd__decap_3 PHY_10107 ();
 sky130_fd_sc_hd__decap_3 PHY_10108 ();
 sky130_fd_sc_hd__decap_3 PHY_10109 ();
 sky130_fd_sc_hd__decap_3 PHY_10110 ();
 sky130_fd_sc_hd__decap_3 PHY_10111 ();
 sky130_fd_sc_hd__decap_3 PHY_10112 ();
 sky130_fd_sc_hd__decap_3 PHY_10113 ();
 sky130_fd_sc_hd__decap_3 PHY_10114 ();
 sky130_fd_sc_hd__decap_3 PHY_10115 ();
 sky130_fd_sc_hd__decap_3 PHY_10116 ();
 sky130_fd_sc_hd__decap_3 PHY_10117 ();
 sky130_fd_sc_hd__decap_3 PHY_10118 ();
 sky130_fd_sc_hd__decap_3 PHY_10119 ();
 sky130_fd_sc_hd__decap_3 PHY_10120 ();
 sky130_fd_sc_hd__decap_3 PHY_10121 ();
 sky130_fd_sc_hd__decap_3 PHY_10122 ();
 sky130_fd_sc_hd__decap_3 PHY_10123 ();
 sky130_fd_sc_hd__decap_3 PHY_10124 ();
 sky130_fd_sc_hd__decap_3 PHY_10125 ();
 sky130_fd_sc_hd__decap_3 PHY_10126 ();
 sky130_fd_sc_hd__decap_3 PHY_10127 ();
 sky130_fd_sc_hd__decap_3 PHY_10128 ();
 sky130_fd_sc_hd__decap_3 PHY_10129 ();
 sky130_fd_sc_hd__decap_3 PHY_10130 ();
 sky130_fd_sc_hd__decap_3 PHY_10131 ();
 sky130_fd_sc_hd__decap_3 PHY_10132 ();
 sky130_fd_sc_hd__decap_3 PHY_10133 ();
 sky130_fd_sc_hd__decap_3 PHY_10134 ();
 sky130_fd_sc_hd__decap_3 PHY_10135 ();
 sky130_fd_sc_hd__decap_3 PHY_10136 ();
 sky130_fd_sc_hd__decap_3 PHY_10137 ();
 sky130_fd_sc_hd__decap_3 PHY_10138 ();
 sky130_fd_sc_hd__decap_3 PHY_10139 ();
 sky130_fd_sc_hd__decap_3 PHY_10140 ();
 sky130_fd_sc_hd__decap_3 PHY_10141 ();
 sky130_fd_sc_hd__decap_3 PHY_10142 ();
 sky130_fd_sc_hd__decap_3 PHY_10143 ();
 sky130_fd_sc_hd__decap_3 PHY_10144 ();
 sky130_fd_sc_hd__decap_3 PHY_10145 ();
 sky130_fd_sc_hd__decap_3 PHY_10146 ();
 sky130_fd_sc_hd__decap_3 PHY_10147 ();
 sky130_fd_sc_hd__decap_3 PHY_10148 ();
 sky130_fd_sc_hd__decap_3 PHY_10149 ();
 sky130_fd_sc_hd__decap_3 PHY_10150 ();
 sky130_fd_sc_hd__decap_3 PHY_10151 ();
 sky130_fd_sc_hd__decap_3 PHY_10152 ();
 sky130_fd_sc_hd__decap_3 PHY_10153 ();
 sky130_fd_sc_hd__decap_3 PHY_10154 ();
 sky130_fd_sc_hd__decap_3 PHY_10155 ();
 sky130_fd_sc_hd__decap_3 PHY_10156 ();
 sky130_fd_sc_hd__decap_3 PHY_10157 ();
 sky130_fd_sc_hd__decap_3 PHY_10158 ();
 sky130_fd_sc_hd__decap_3 PHY_10159 ();
 sky130_fd_sc_hd__decap_3 PHY_10160 ();
 sky130_fd_sc_hd__decap_3 PHY_10161 ();
 sky130_fd_sc_hd__decap_3 PHY_10162 ();
 sky130_fd_sc_hd__decap_3 PHY_10163 ();
 sky130_fd_sc_hd__decap_3 PHY_10164 ();
 sky130_fd_sc_hd__decap_3 PHY_10165 ();
 sky130_fd_sc_hd__decap_3 PHY_10166 ();
 sky130_fd_sc_hd__decap_3 PHY_10167 ();
 sky130_fd_sc_hd__decap_3 PHY_10168 ();
 sky130_fd_sc_hd__decap_3 PHY_10169 ();
 sky130_fd_sc_hd__decap_3 PHY_10170 ();
 sky130_fd_sc_hd__decap_3 PHY_10171 ();
 sky130_fd_sc_hd__decap_3 PHY_10172 ();
 sky130_fd_sc_hd__decap_3 PHY_10173 ();
 sky130_fd_sc_hd__decap_3 PHY_10174 ();
 sky130_fd_sc_hd__decap_3 PHY_10175 ();
 sky130_fd_sc_hd__decap_3 PHY_10176 ();
 sky130_fd_sc_hd__decap_3 PHY_10177 ();
 sky130_fd_sc_hd__decap_3 PHY_10178 ();
 sky130_fd_sc_hd__decap_3 PHY_10179 ();
 sky130_fd_sc_hd__decap_3 PHY_10180 ();
 sky130_fd_sc_hd__decap_3 PHY_10181 ();
 sky130_fd_sc_hd__decap_3 PHY_10182 ();
 sky130_fd_sc_hd__decap_3 PHY_10183 ();
 sky130_fd_sc_hd__decap_3 PHY_10184 ();
 sky130_fd_sc_hd__decap_3 PHY_10185 ();
 sky130_fd_sc_hd__decap_3 PHY_10186 ();
 sky130_fd_sc_hd__decap_3 PHY_10187 ();
 sky130_fd_sc_hd__decap_3 PHY_10188 ();
 sky130_fd_sc_hd__decap_3 PHY_10189 ();
 sky130_fd_sc_hd__decap_3 PHY_10190 ();
 sky130_fd_sc_hd__decap_3 PHY_10191 ();
 sky130_fd_sc_hd__decap_3 PHY_10192 ();
 sky130_fd_sc_hd__decap_3 PHY_10193 ();
 sky130_fd_sc_hd__decap_3 PHY_10194 ();
 sky130_fd_sc_hd__decap_3 PHY_10195 ();
 sky130_fd_sc_hd__decap_3 PHY_10196 ();
 sky130_fd_sc_hd__decap_3 PHY_10197 ();
 sky130_fd_sc_hd__decap_3 PHY_10198 ();
 sky130_fd_sc_hd__decap_3 PHY_10199 ();
 sky130_fd_sc_hd__decap_3 PHY_10200 ();
 sky130_fd_sc_hd__decap_3 PHY_10201 ();
 sky130_fd_sc_hd__decap_3 PHY_10202 ();
 sky130_fd_sc_hd__decap_3 PHY_10203 ();
 sky130_fd_sc_hd__decap_3 PHY_10204 ();
 sky130_fd_sc_hd__decap_3 PHY_10205 ();
 sky130_fd_sc_hd__decap_3 PHY_10206 ();
 sky130_fd_sc_hd__decap_3 PHY_10207 ();
 sky130_fd_sc_hd__decap_3 PHY_10208 ();
 sky130_fd_sc_hd__decap_3 PHY_10209 ();
 sky130_fd_sc_hd__decap_3 PHY_10210 ();
 sky130_fd_sc_hd__decap_3 PHY_10211 ();
 sky130_fd_sc_hd__decap_3 PHY_10212 ();
 sky130_fd_sc_hd__decap_3 PHY_10213 ();
 sky130_fd_sc_hd__decap_3 PHY_10214 ();
 sky130_fd_sc_hd__decap_3 PHY_10215 ();
 sky130_fd_sc_hd__decap_3 PHY_10216 ();
 sky130_fd_sc_hd__decap_3 PHY_10217 ();
 sky130_fd_sc_hd__decap_3 PHY_10218 ();
 sky130_fd_sc_hd__decap_3 PHY_10219 ();
 sky130_fd_sc_hd__decap_3 PHY_10220 ();
 sky130_fd_sc_hd__decap_3 PHY_10221 ();
 sky130_fd_sc_hd__decap_3 PHY_10222 ();
 sky130_fd_sc_hd__decap_3 PHY_10223 ();
 sky130_fd_sc_hd__decap_3 PHY_10224 ();
 sky130_fd_sc_hd__decap_3 PHY_10225 ();
 sky130_fd_sc_hd__decap_3 PHY_10226 ();
 sky130_fd_sc_hd__decap_3 PHY_10227 ();
 sky130_fd_sc_hd__decap_3 PHY_10228 ();
 sky130_fd_sc_hd__decap_3 PHY_10229 ();
 sky130_fd_sc_hd__decap_3 PHY_10230 ();
 sky130_fd_sc_hd__decap_3 PHY_10231 ();
 sky130_fd_sc_hd__decap_3 PHY_10232 ();
 sky130_fd_sc_hd__decap_3 PHY_10233 ();
 sky130_fd_sc_hd__decap_3 PHY_10234 ();
 sky130_fd_sc_hd__decap_3 PHY_10235 ();
 sky130_fd_sc_hd__decap_3 PHY_10236 ();
 sky130_fd_sc_hd__decap_3 PHY_10237 ();
 sky130_fd_sc_hd__decap_3 PHY_10238 ();
 sky130_fd_sc_hd__decap_3 PHY_10239 ();
 sky130_fd_sc_hd__decap_3 PHY_10240 ();
 sky130_fd_sc_hd__decap_3 PHY_10241 ();
 sky130_fd_sc_hd__decap_3 PHY_10242 ();
 sky130_fd_sc_hd__decap_3 PHY_10243 ();
 sky130_fd_sc_hd__decap_3 PHY_10244 ();
 sky130_fd_sc_hd__decap_3 PHY_10245 ();
 sky130_fd_sc_hd__decap_3 PHY_10246 ();
 sky130_fd_sc_hd__decap_3 PHY_10247 ();
 sky130_fd_sc_hd__decap_3 PHY_10248 ();
 sky130_fd_sc_hd__decap_3 PHY_10249 ();
 sky130_fd_sc_hd__decap_3 PHY_10250 ();
 sky130_fd_sc_hd__decap_3 PHY_10251 ();
 sky130_fd_sc_hd__decap_3 PHY_10252 ();
 sky130_fd_sc_hd__decap_3 PHY_10253 ();
 sky130_fd_sc_hd__decap_3 PHY_10254 ();
 sky130_fd_sc_hd__decap_3 PHY_10255 ();
 sky130_fd_sc_hd__decap_3 PHY_10256 ();
 sky130_fd_sc_hd__decap_3 PHY_10257 ();
 sky130_fd_sc_hd__decap_3 PHY_10258 ();
 sky130_fd_sc_hd__decap_3 PHY_10259 ();
 sky130_fd_sc_hd__decap_3 PHY_10260 ();
 sky130_fd_sc_hd__decap_3 PHY_10261 ();
 sky130_fd_sc_hd__decap_3 PHY_10262 ();
 sky130_fd_sc_hd__decap_3 PHY_10263 ();
 sky130_fd_sc_hd__decap_3 PHY_10264 ();
 sky130_fd_sc_hd__decap_3 PHY_10265 ();
 sky130_fd_sc_hd__decap_3 PHY_10266 ();
 sky130_fd_sc_hd__decap_3 PHY_10267 ();
 sky130_fd_sc_hd__decap_3 PHY_10268 ();
 sky130_fd_sc_hd__decap_3 PHY_10269 ();
 sky130_fd_sc_hd__decap_3 PHY_10270 ();
 sky130_fd_sc_hd__decap_3 PHY_10271 ();
 sky130_fd_sc_hd__decap_3 PHY_10272 ();
 sky130_fd_sc_hd__decap_3 PHY_10273 ();
 sky130_fd_sc_hd__decap_3 PHY_10274 ();
 sky130_fd_sc_hd__decap_3 PHY_10275 ();
 sky130_fd_sc_hd__decap_3 PHY_10276 ();
 sky130_fd_sc_hd__decap_3 PHY_10277 ();
 sky130_fd_sc_hd__decap_3 PHY_10278 ();
 sky130_fd_sc_hd__decap_3 PHY_10279 ();
 sky130_fd_sc_hd__decap_3 PHY_10280 ();
 sky130_fd_sc_hd__decap_3 PHY_10281 ();
 sky130_fd_sc_hd__decap_3 PHY_10282 ();
 sky130_fd_sc_hd__decap_3 PHY_10283 ();
 sky130_fd_sc_hd__decap_3 PHY_10284 ();
 sky130_fd_sc_hd__decap_3 PHY_10285 ();
 sky130_fd_sc_hd__decap_3 PHY_10286 ();
 sky130_fd_sc_hd__decap_3 PHY_10287 ();
 sky130_fd_sc_hd__decap_3 PHY_10288 ();
 sky130_fd_sc_hd__decap_3 PHY_10289 ();
 sky130_fd_sc_hd__decap_3 PHY_10290 ();
 sky130_fd_sc_hd__decap_3 PHY_10291 ();
 sky130_fd_sc_hd__decap_3 PHY_10292 ();
 sky130_fd_sc_hd__decap_3 PHY_10293 ();
 sky130_fd_sc_hd__decap_3 PHY_10294 ();
 sky130_fd_sc_hd__decap_3 PHY_10295 ();
 sky130_fd_sc_hd__decap_3 PHY_10296 ();
 sky130_fd_sc_hd__decap_3 PHY_10297 ();
 sky130_fd_sc_hd__decap_3 PHY_10298 ();
 sky130_fd_sc_hd__decap_3 PHY_10299 ();
 sky130_fd_sc_hd__decap_3 PHY_10300 ();
 sky130_fd_sc_hd__decap_3 PHY_10301 ();
 sky130_fd_sc_hd__decap_3 PHY_10302 ();
 sky130_fd_sc_hd__decap_3 PHY_10303 ();
 sky130_fd_sc_hd__decap_3 PHY_10304 ();
 sky130_fd_sc_hd__decap_3 PHY_10305 ();
 sky130_fd_sc_hd__decap_3 PHY_10306 ();
 sky130_fd_sc_hd__decap_3 PHY_10307 ();
 sky130_fd_sc_hd__decap_3 PHY_10308 ();
 sky130_fd_sc_hd__decap_3 PHY_10309 ();
 sky130_fd_sc_hd__decap_3 PHY_10310 ();
 sky130_fd_sc_hd__decap_3 PHY_10311 ();
 sky130_fd_sc_hd__decap_3 PHY_10312 ();
 sky130_fd_sc_hd__decap_3 PHY_10313 ();
 sky130_fd_sc_hd__decap_3 PHY_10314 ();
 sky130_fd_sc_hd__decap_3 PHY_10315 ();
 sky130_fd_sc_hd__decap_3 PHY_10316 ();
 sky130_fd_sc_hd__decap_3 PHY_10317 ();
 sky130_fd_sc_hd__decap_3 PHY_10318 ();
 sky130_fd_sc_hd__decap_3 PHY_10319 ();
 sky130_fd_sc_hd__decap_3 PHY_10320 ();
 sky130_fd_sc_hd__decap_3 PHY_10321 ();
 sky130_fd_sc_hd__decap_3 PHY_10322 ();
 sky130_fd_sc_hd__decap_3 PHY_10323 ();
 sky130_fd_sc_hd__decap_3 PHY_10324 ();
 sky130_fd_sc_hd__decap_3 PHY_10325 ();
 sky130_fd_sc_hd__decap_3 PHY_10326 ();
 sky130_fd_sc_hd__decap_3 PHY_10327 ();
 sky130_fd_sc_hd__decap_3 PHY_10328 ();
 sky130_fd_sc_hd__decap_3 PHY_10329 ();
 sky130_fd_sc_hd__decap_3 PHY_10330 ();
 sky130_fd_sc_hd__decap_3 PHY_10331 ();
 sky130_fd_sc_hd__decap_3 PHY_10332 ();
 sky130_fd_sc_hd__decap_3 PHY_10333 ();
 sky130_fd_sc_hd__decap_3 PHY_10334 ();
 sky130_fd_sc_hd__decap_3 PHY_10335 ();
 sky130_fd_sc_hd__decap_3 PHY_10336 ();
 sky130_fd_sc_hd__decap_3 PHY_10337 ();
 sky130_fd_sc_hd__decap_3 PHY_10338 ();
 sky130_fd_sc_hd__decap_3 PHY_10339 ();
 sky130_fd_sc_hd__decap_3 PHY_10340 ();
 sky130_fd_sc_hd__decap_3 PHY_10341 ();
 sky130_fd_sc_hd__decap_3 PHY_10342 ();
 sky130_fd_sc_hd__decap_3 PHY_10343 ();
 sky130_fd_sc_hd__decap_3 PHY_10344 ();
 sky130_fd_sc_hd__decap_3 PHY_10345 ();
 sky130_fd_sc_hd__decap_3 PHY_10346 ();
 sky130_fd_sc_hd__decap_3 PHY_10347 ();
 sky130_fd_sc_hd__decap_3 PHY_10348 ();
 sky130_fd_sc_hd__decap_3 PHY_10349 ();
 sky130_fd_sc_hd__decap_3 PHY_10350 ();
 sky130_fd_sc_hd__decap_3 PHY_10351 ();
 sky130_fd_sc_hd__decap_3 PHY_10352 ();
 sky130_fd_sc_hd__decap_3 PHY_10353 ();
 sky130_fd_sc_hd__decap_3 PHY_10354 ();
 sky130_fd_sc_hd__decap_3 PHY_10355 ();
 sky130_fd_sc_hd__decap_3 PHY_10356 ();
 sky130_fd_sc_hd__decap_3 PHY_10357 ();
 sky130_fd_sc_hd__decap_3 PHY_10358 ();
 sky130_fd_sc_hd__decap_3 PHY_10359 ();
 sky130_fd_sc_hd__decap_3 PHY_10360 ();
 sky130_fd_sc_hd__decap_3 PHY_10361 ();
 sky130_fd_sc_hd__decap_3 PHY_10362 ();
 sky130_fd_sc_hd__decap_3 PHY_10363 ();
 sky130_fd_sc_hd__decap_3 PHY_10364 ();
 sky130_fd_sc_hd__decap_3 PHY_10365 ();
 sky130_fd_sc_hd__decap_3 PHY_10366 ();
 sky130_fd_sc_hd__decap_3 PHY_10367 ();
 sky130_fd_sc_hd__decap_3 PHY_10368 ();
 sky130_fd_sc_hd__decap_3 PHY_10369 ();
 sky130_fd_sc_hd__decap_3 PHY_10370 ();
 sky130_fd_sc_hd__decap_3 PHY_10371 ();
 sky130_fd_sc_hd__decap_3 PHY_10372 ();
 sky130_fd_sc_hd__decap_3 PHY_10373 ();
 sky130_fd_sc_hd__decap_3 PHY_10374 ();
 sky130_fd_sc_hd__decap_3 PHY_10375 ();
 sky130_fd_sc_hd__decap_3 PHY_10376 ();
 sky130_fd_sc_hd__decap_3 PHY_10377 ();
 sky130_fd_sc_hd__decap_3 PHY_10378 ();
 sky130_fd_sc_hd__decap_3 PHY_10379 ();
 sky130_fd_sc_hd__decap_3 PHY_10380 ();
 sky130_fd_sc_hd__decap_3 PHY_10381 ();
 sky130_fd_sc_hd__decap_3 PHY_10382 ();
 sky130_fd_sc_hd__decap_3 PHY_10383 ();
 sky130_fd_sc_hd__decap_3 PHY_10384 ();
 sky130_fd_sc_hd__decap_3 PHY_10385 ();
 sky130_fd_sc_hd__decap_3 PHY_10386 ();
 sky130_fd_sc_hd__decap_3 PHY_10387 ();
 sky130_fd_sc_hd__decap_3 PHY_10388 ();
 sky130_fd_sc_hd__decap_3 PHY_10389 ();
 sky130_fd_sc_hd__decap_3 PHY_10390 ();
 sky130_fd_sc_hd__decap_3 PHY_10391 ();
 sky130_fd_sc_hd__decap_3 PHY_10392 ();
 sky130_fd_sc_hd__decap_3 PHY_10393 ();
 sky130_fd_sc_hd__decap_3 PHY_10394 ();
 sky130_fd_sc_hd__decap_3 PHY_10395 ();
 sky130_fd_sc_hd__decap_3 PHY_10396 ();
 sky130_fd_sc_hd__decap_3 PHY_10397 ();
 sky130_fd_sc_hd__decap_3 PHY_10398 ();
 sky130_fd_sc_hd__decap_3 PHY_10399 ();
 sky130_fd_sc_hd__decap_3 PHY_10400 ();
 sky130_fd_sc_hd__decap_3 PHY_10401 ();
 sky130_fd_sc_hd__decap_3 PHY_10402 ();
 sky130_fd_sc_hd__decap_3 PHY_10403 ();
 sky130_fd_sc_hd__decap_3 PHY_10404 ();
 sky130_fd_sc_hd__decap_3 PHY_10405 ();
 sky130_fd_sc_hd__decap_3 PHY_10406 ();
 sky130_fd_sc_hd__decap_3 PHY_10407 ();
 sky130_fd_sc_hd__decap_3 PHY_10408 ();
 sky130_fd_sc_hd__decap_3 PHY_10409 ();
 sky130_fd_sc_hd__decap_3 PHY_10410 ();
 sky130_fd_sc_hd__decap_3 PHY_10411 ();
 sky130_fd_sc_hd__decap_3 PHY_10412 ();
 sky130_fd_sc_hd__decap_3 PHY_10413 ();
 sky130_fd_sc_hd__decap_3 PHY_10414 ();
 sky130_fd_sc_hd__decap_3 PHY_10415 ();
 sky130_fd_sc_hd__decap_3 PHY_10416 ();
 sky130_fd_sc_hd__decap_3 PHY_10417 ();
 sky130_fd_sc_hd__decap_3 PHY_10418 ();
 sky130_fd_sc_hd__decap_3 PHY_10419 ();
 sky130_fd_sc_hd__decap_3 PHY_10420 ();
 sky130_fd_sc_hd__decap_3 PHY_10421 ();
 sky130_fd_sc_hd__decap_3 PHY_10422 ();
 sky130_fd_sc_hd__decap_3 PHY_10423 ();
 sky130_fd_sc_hd__decap_3 PHY_10424 ();
 sky130_fd_sc_hd__decap_3 PHY_10425 ();
 sky130_fd_sc_hd__decap_3 PHY_10426 ();
 sky130_fd_sc_hd__decap_3 PHY_10427 ();
 sky130_fd_sc_hd__decap_3 PHY_10428 ();
 sky130_fd_sc_hd__decap_3 PHY_10429 ();
 sky130_fd_sc_hd__decap_3 PHY_10430 ();
 sky130_fd_sc_hd__decap_3 PHY_10431 ();
 sky130_fd_sc_hd__decap_3 PHY_10432 ();
 sky130_fd_sc_hd__decap_3 PHY_10433 ();
 sky130_fd_sc_hd__decap_3 PHY_10434 ();
 sky130_fd_sc_hd__decap_3 PHY_10435 ();
 sky130_fd_sc_hd__decap_3 PHY_10436 ();
 sky130_fd_sc_hd__decap_3 PHY_10437 ();
 sky130_fd_sc_hd__decap_3 PHY_10438 ();
 sky130_fd_sc_hd__decap_3 PHY_10439 ();
 sky130_fd_sc_hd__decap_3 PHY_10440 ();
 sky130_fd_sc_hd__decap_3 PHY_10441 ();
 sky130_fd_sc_hd__decap_3 PHY_10442 ();
 sky130_fd_sc_hd__decap_3 PHY_10443 ();
 sky130_fd_sc_hd__decap_3 PHY_10444 ();
 sky130_fd_sc_hd__decap_3 PHY_10445 ();
 sky130_fd_sc_hd__decap_3 PHY_10446 ();
 sky130_fd_sc_hd__decap_3 PHY_10447 ();
 sky130_fd_sc_hd__decap_3 PHY_10448 ();
 sky130_fd_sc_hd__decap_3 PHY_10449 ();
 sky130_fd_sc_hd__decap_3 PHY_10450 ();
 sky130_fd_sc_hd__decap_3 PHY_10451 ();
 sky130_fd_sc_hd__decap_3 PHY_10452 ();
 sky130_fd_sc_hd__decap_3 PHY_10453 ();
 sky130_fd_sc_hd__decap_3 PHY_10454 ();
 sky130_fd_sc_hd__decap_3 PHY_10455 ();
 sky130_fd_sc_hd__decap_3 PHY_10456 ();
 sky130_fd_sc_hd__decap_3 PHY_10457 ();
 sky130_fd_sc_hd__decap_3 PHY_10458 ();
 sky130_fd_sc_hd__decap_3 PHY_10459 ();
 sky130_fd_sc_hd__decap_3 PHY_10460 ();
 sky130_fd_sc_hd__decap_3 PHY_10461 ();
 sky130_fd_sc_hd__decap_3 PHY_10462 ();
 sky130_fd_sc_hd__decap_3 PHY_10463 ();
 sky130_fd_sc_hd__decap_3 PHY_10464 ();
 sky130_fd_sc_hd__decap_3 PHY_10465 ();
 sky130_fd_sc_hd__decap_3 PHY_10466 ();
 sky130_fd_sc_hd__decap_3 PHY_10467 ();
 sky130_fd_sc_hd__decap_3 PHY_10468 ();
 sky130_fd_sc_hd__decap_3 PHY_10469 ();
 sky130_fd_sc_hd__decap_3 PHY_10470 ();
 sky130_fd_sc_hd__decap_3 PHY_10471 ();
 sky130_fd_sc_hd__decap_3 PHY_10472 ();
 sky130_fd_sc_hd__decap_3 PHY_10473 ();
 sky130_fd_sc_hd__decap_3 PHY_10474 ();
 sky130_fd_sc_hd__decap_3 PHY_10475 ();
 sky130_fd_sc_hd__decap_3 PHY_10476 ();
 sky130_fd_sc_hd__decap_3 PHY_10477 ();
 sky130_fd_sc_hd__decap_3 PHY_10478 ();
 sky130_fd_sc_hd__decap_3 PHY_10479 ();
 sky130_fd_sc_hd__decap_3 PHY_10480 ();
 sky130_fd_sc_hd__decap_3 PHY_10481 ();
 sky130_fd_sc_hd__decap_3 PHY_10482 ();
 sky130_fd_sc_hd__decap_3 PHY_10483 ();
 sky130_fd_sc_hd__decap_3 PHY_10484 ();
 sky130_fd_sc_hd__decap_3 PHY_10485 ();
 sky130_fd_sc_hd__decap_3 PHY_10486 ();
 sky130_fd_sc_hd__decap_3 PHY_10487 ();
 sky130_fd_sc_hd__decap_3 PHY_10488 ();
 sky130_fd_sc_hd__decap_3 PHY_10489 ();
 sky130_fd_sc_hd__decap_3 PHY_10490 ();
 sky130_fd_sc_hd__decap_3 PHY_10491 ();
 sky130_fd_sc_hd__decap_3 PHY_10492 ();
 sky130_fd_sc_hd__decap_3 PHY_10493 ();
 sky130_fd_sc_hd__decap_3 PHY_10494 ();
 sky130_fd_sc_hd__decap_3 PHY_10495 ();
 sky130_fd_sc_hd__decap_3 PHY_10496 ();
 sky130_fd_sc_hd__decap_3 PHY_10497 ();
 sky130_fd_sc_hd__decap_3 PHY_10498 ();
 sky130_fd_sc_hd__decap_3 PHY_10499 ();
 sky130_fd_sc_hd__decap_3 PHY_10500 ();
 sky130_fd_sc_hd__decap_3 PHY_10501 ();
 sky130_fd_sc_hd__decap_3 PHY_10502 ();
 sky130_fd_sc_hd__decap_3 PHY_10503 ();
 sky130_fd_sc_hd__decap_3 PHY_10504 ();
 sky130_fd_sc_hd__decap_3 PHY_10505 ();
 sky130_fd_sc_hd__decap_3 PHY_10506 ();
 sky130_fd_sc_hd__decap_3 PHY_10507 ();
 sky130_fd_sc_hd__decap_3 PHY_10508 ();
 sky130_fd_sc_hd__decap_3 PHY_10509 ();
 sky130_fd_sc_hd__decap_3 PHY_10510 ();
 sky130_fd_sc_hd__decap_3 PHY_10511 ();
 sky130_fd_sc_hd__decap_3 PHY_10512 ();
 sky130_fd_sc_hd__decap_3 PHY_10513 ();
 sky130_fd_sc_hd__decap_3 PHY_10514 ();
 sky130_fd_sc_hd__decap_3 PHY_10515 ();
 sky130_fd_sc_hd__decap_3 PHY_10516 ();
 sky130_fd_sc_hd__decap_3 PHY_10517 ();
 sky130_fd_sc_hd__decap_3 PHY_10518 ();
 sky130_fd_sc_hd__decap_3 PHY_10519 ();
 sky130_fd_sc_hd__decap_3 PHY_10520 ();
 sky130_fd_sc_hd__decap_3 PHY_10521 ();
 sky130_fd_sc_hd__decap_3 PHY_10522 ();
 sky130_fd_sc_hd__decap_3 PHY_10523 ();
 sky130_fd_sc_hd__decap_3 PHY_10524 ();
 sky130_fd_sc_hd__decap_3 PHY_10525 ();
 sky130_fd_sc_hd__decap_3 PHY_10526 ();
 sky130_fd_sc_hd__decap_3 PHY_10527 ();
 sky130_fd_sc_hd__decap_3 PHY_10528 ();
 sky130_fd_sc_hd__decap_3 PHY_10529 ();
 sky130_fd_sc_hd__decap_3 PHY_10530 ();
 sky130_fd_sc_hd__decap_3 PHY_10531 ();
 sky130_fd_sc_hd__decap_3 PHY_10532 ();
 sky130_fd_sc_hd__decap_3 PHY_10533 ();
 sky130_fd_sc_hd__decap_3 PHY_10534 ();
 sky130_fd_sc_hd__decap_3 PHY_10535 ();
 sky130_fd_sc_hd__decap_3 PHY_10536 ();
 sky130_fd_sc_hd__decap_3 PHY_10537 ();
 sky130_fd_sc_hd__decap_3 PHY_10538 ();
 sky130_fd_sc_hd__decap_3 PHY_10539 ();
 sky130_fd_sc_hd__decap_3 PHY_10540 ();
 sky130_fd_sc_hd__decap_3 PHY_10541 ();
 sky130_fd_sc_hd__decap_3 PHY_10542 ();
 sky130_fd_sc_hd__decap_3 PHY_10543 ();
 sky130_fd_sc_hd__decap_3 PHY_10544 ();
 sky130_fd_sc_hd__decap_3 PHY_10545 ();
 sky130_fd_sc_hd__decap_3 PHY_10546 ();
 sky130_fd_sc_hd__decap_3 PHY_10547 ();
 sky130_fd_sc_hd__decap_3 PHY_10548 ();
 sky130_fd_sc_hd__decap_3 PHY_10549 ();
 sky130_fd_sc_hd__decap_3 PHY_10550 ();
 sky130_fd_sc_hd__decap_3 PHY_10551 ();
 sky130_fd_sc_hd__decap_3 PHY_10552 ();
 sky130_fd_sc_hd__decap_3 PHY_10553 ();
 sky130_fd_sc_hd__decap_3 PHY_10554 ();
 sky130_fd_sc_hd__decap_3 PHY_10555 ();
 sky130_fd_sc_hd__decap_3 PHY_10556 ();
 sky130_fd_sc_hd__decap_3 PHY_10557 ();
 sky130_fd_sc_hd__decap_3 PHY_10558 ();
 sky130_fd_sc_hd__decap_3 PHY_10559 ();
 sky130_fd_sc_hd__decap_3 PHY_10560 ();
 sky130_fd_sc_hd__decap_3 PHY_10561 ();
 sky130_fd_sc_hd__decap_3 PHY_10562 ();
 sky130_fd_sc_hd__decap_3 PHY_10563 ();
 sky130_fd_sc_hd__decap_3 PHY_10564 ();
 sky130_fd_sc_hd__decap_3 PHY_10565 ();
 sky130_fd_sc_hd__decap_3 PHY_10566 ();
 sky130_fd_sc_hd__decap_3 PHY_10567 ();
 sky130_fd_sc_hd__decap_3 PHY_10568 ();
 sky130_fd_sc_hd__decap_3 PHY_10569 ();
 sky130_fd_sc_hd__decap_3 PHY_10570 ();
 sky130_fd_sc_hd__decap_3 PHY_10571 ();
 sky130_fd_sc_hd__decap_3 PHY_10572 ();
 sky130_fd_sc_hd__decap_3 PHY_10573 ();
 sky130_fd_sc_hd__decap_3 PHY_10574 ();
 sky130_fd_sc_hd__decap_3 PHY_10575 ();
 sky130_fd_sc_hd__decap_3 PHY_10576 ();
 sky130_fd_sc_hd__decap_3 PHY_10577 ();
 sky130_fd_sc_hd__decap_3 PHY_10578 ();
 sky130_fd_sc_hd__decap_3 PHY_10579 ();
 sky130_fd_sc_hd__decap_3 PHY_10580 ();
 sky130_fd_sc_hd__decap_3 PHY_10581 ();
 sky130_fd_sc_hd__decap_3 PHY_10582 ();
 sky130_fd_sc_hd__decap_3 PHY_10583 ();
 sky130_fd_sc_hd__decap_3 PHY_10584 ();
 sky130_fd_sc_hd__decap_3 PHY_10585 ();
 sky130_fd_sc_hd__decap_3 PHY_10586 ();
 sky130_fd_sc_hd__decap_3 PHY_10587 ();
 sky130_fd_sc_hd__decap_3 PHY_10588 ();
 sky130_fd_sc_hd__decap_3 PHY_10589 ();
 sky130_fd_sc_hd__decap_3 PHY_10590 ();
 sky130_fd_sc_hd__decap_3 PHY_10591 ();
 sky130_fd_sc_hd__decap_3 PHY_10592 ();
 sky130_fd_sc_hd__decap_3 PHY_10593 ();
 sky130_fd_sc_hd__decap_3 PHY_10594 ();
 sky130_fd_sc_hd__decap_3 PHY_10595 ();
 sky130_fd_sc_hd__decap_3 PHY_10596 ();
 sky130_fd_sc_hd__decap_3 PHY_10597 ();
 sky130_fd_sc_hd__decap_3 PHY_10598 ();
 sky130_fd_sc_hd__decap_3 PHY_10599 ();
 sky130_fd_sc_hd__decap_3 PHY_10600 ();
 sky130_fd_sc_hd__decap_3 PHY_10601 ();
 sky130_fd_sc_hd__decap_3 PHY_10602 ();
 sky130_fd_sc_hd__decap_3 PHY_10603 ();
 sky130_fd_sc_hd__decap_3 PHY_10604 ();
 sky130_fd_sc_hd__decap_3 PHY_10605 ();
 sky130_fd_sc_hd__decap_3 PHY_10606 ();
 sky130_fd_sc_hd__decap_3 PHY_10607 ();
 sky130_fd_sc_hd__decap_3 PHY_10608 ();
 sky130_fd_sc_hd__decap_3 PHY_10609 ();
 sky130_fd_sc_hd__decap_3 PHY_10610 ();
 sky130_fd_sc_hd__decap_3 PHY_10611 ();
 sky130_fd_sc_hd__decap_3 PHY_10612 ();
 sky130_fd_sc_hd__decap_3 PHY_10613 ();
 sky130_fd_sc_hd__decap_3 PHY_10614 ();
 sky130_fd_sc_hd__decap_3 PHY_10615 ();
 sky130_fd_sc_hd__decap_3 PHY_10616 ();
 sky130_fd_sc_hd__decap_3 PHY_10617 ();
 sky130_fd_sc_hd__decap_3 PHY_10618 ();
 sky130_fd_sc_hd__decap_3 PHY_10619 ();
 sky130_fd_sc_hd__decap_3 PHY_10620 ();
 sky130_fd_sc_hd__decap_3 PHY_10621 ();
 sky130_fd_sc_hd__decap_3 PHY_10622 ();
 sky130_fd_sc_hd__decap_3 PHY_10623 ();
 sky130_fd_sc_hd__decap_3 PHY_10624 ();
 sky130_fd_sc_hd__decap_3 PHY_10625 ();
 sky130_fd_sc_hd__decap_3 PHY_10626 ();
 sky130_fd_sc_hd__decap_3 PHY_10627 ();
 sky130_fd_sc_hd__decap_3 PHY_10628 ();
 sky130_fd_sc_hd__decap_3 PHY_10629 ();
 sky130_fd_sc_hd__decap_3 PHY_10630 ();
 sky130_fd_sc_hd__decap_3 PHY_10631 ();
 sky130_fd_sc_hd__decap_3 PHY_10632 ();
 sky130_fd_sc_hd__decap_3 PHY_10633 ();
 sky130_fd_sc_hd__decap_3 PHY_10634 ();
 sky130_fd_sc_hd__decap_3 PHY_10635 ();
 sky130_fd_sc_hd__decap_3 PHY_10636 ();
 sky130_fd_sc_hd__decap_3 PHY_10637 ();
 sky130_fd_sc_hd__decap_3 PHY_10638 ();
 sky130_fd_sc_hd__decap_3 PHY_10639 ();
 sky130_fd_sc_hd__decap_3 PHY_10640 ();
 sky130_fd_sc_hd__decap_3 PHY_10641 ();
 sky130_fd_sc_hd__decap_3 PHY_10642 ();
 sky130_fd_sc_hd__decap_3 PHY_10643 ();
 sky130_fd_sc_hd__decap_3 PHY_10644 ();
 sky130_fd_sc_hd__decap_3 PHY_10645 ();
 sky130_fd_sc_hd__decap_3 PHY_10646 ();
 sky130_fd_sc_hd__decap_3 PHY_10647 ();
 sky130_fd_sc_hd__decap_3 PHY_10648 ();
 sky130_fd_sc_hd__decap_3 PHY_10649 ();
 sky130_fd_sc_hd__decap_3 PHY_10650 ();
 sky130_fd_sc_hd__decap_3 PHY_10651 ();
 sky130_fd_sc_hd__decap_3 PHY_10652 ();
 sky130_fd_sc_hd__decap_3 PHY_10653 ();
 sky130_fd_sc_hd__decap_3 PHY_10654 ();
 sky130_fd_sc_hd__decap_3 PHY_10655 ();
 sky130_fd_sc_hd__decap_3 PHY_10656 ();
 sky130_fd_sc_hd__decap_3 PHY_10657 ();
 sky130_fd_sc_hd__decap_3 PHY_10658 ();
 sky130_fd_sc_hd__decap_3 PHY_10659 ();
 sky130_fd_sc_hd__decap_3 PHY_10660 ();
 sky130_fd_sc_hd__decap_3 PHY_10661 ();
 sky130_fd_sc_hd__decap_3 PHY_10662 ();
 sky130_fd_sc_hd__decap_3 PHY_10663 ();
 sky130_fd_sc_hd__decap_3 PHY_10664 ();
 sky130_fd_sc_hd__decap_3 PHY_10665 ();
 sky130_fd_sc_hd__decap_3 PHY_10666 ();
 sky130_fd_sc_hd__decap_3 PHY_10667 ();
 sky130_fd_sc_hd__decap_3 PHY_10668 ();
 sky130_fd_sc_hd__decap_3 PHY_10669 ();
 sky130_fd_sc_hd__decap_3 PHY_10670 ();
 sky130_fd_sc_hd__decap_3 PHY_10671 ();
 sky130_fd_sc_hd__decap_3 PHY_10672 ();
 sky130_fd_sc_hd__decap_3 PHY_10673 ();
 sky130_fd_sc_hd__decap_3 PHY_10674 ();
 sky130_fd_sc_hd__decap_3 PHY_10675 ();
 sky130_fd_sc_hd__decap_3 PHY_10676 ();
 sky130_fd_sc_hd__decap_3 PHY_10677 ();
 sky130_fd_sc_hd__decap_3 PHY_10678 ();
 sky130_fd_sc_hd__decap_3 PHY_10679 ();
 sky130_fd_sc_hd__decap_3 PHY_10680 ();
 sky130_fd_sc_hd__decap_3 PHY_10681 ();
 sky130_fd_sc_hd__decap_3 PHY_10682 ();
 sky130_fd_sc_hd__decap_3 PHY_10683 ();
 sky130_fd_sc_hd__decap_3 PHY_10684 ();
 sky130_fd_sc_hd__decap_3 PHY_10685 ();
 sky130_fd_sc_hd__decap_3 PHY_10686 ();
 sky130_fd_sc_hd__decap_3 PHY_10687 ();
 sky130_fd_sc_hd__decap_3 PHY_10688 ();
 sky130_fd_sc_hd__decap_3 PHY_10689 ();
 sky130_fd_sc_hd__decap_3 PHY_10690 ();
 sky130_fd_sc_hd__decap_3 PHY_10691 ();
 sky130_fd_sc_hd__decap_3 PHY_10692 ();
 sky130_fd_sc_hd__decap_3 PHY_10693 ();
 sky130_fd_sc_hd__decap_3 PHY_10694 ();
 sky130_fd_sc_hd__decap_3 PHY_10695 ();
 sky130_fd_sc_hd__decap_3 PHY_10696 ();
 sky130_fd_sc_hd__decap_3 PHY_10697 ();
 sky130_fd_sc_hd__decap_3 PHY_10698 ();
 sky130_fd_sc_hd__decap_3 PHY_10699 ();
 sky130_fd_sc_hd__decap_3 PHY_10700 ();
 sky130_fd_sc_hd__decap_3 PHY_10701 ();
 sky130_fd_sc_hd__decap_3 PHY_10702 ();
 sky130_fd_sc_hd__decap_3 PHY_10703 ();
 sky130_fd_sc_hd__decap_3 PHY_10704 ();
 sky130_fd_sc_hd__decap_3 PHY_10705 ();
 sky130_fd_sc_hd__decap_3 PHY_10706 ();
 sky130_fd_sc_hd__decap_3 PHY_10707 ();
 sky130_fd_sc_hd__decap_3 PHY_10708 ();
 sky130_fd_sc_hd__decap_3 PHY_10709 ();
 sky130_fd_sc_hd__decap_3 PHY_10710 ();
 sky130_fd_sc_hd__decap_3 PHY_10711 ();
 sky130_fd_sc_hd__decap_3 PHY_10712 ();
 sky130_fd_sc_hd__decap_3 PHY_10713 ();
 sky130_fd_sc_hd__decap_3 PHY_10714 ();
 sky130_fd_sc_hd__decap_3 PHY_10715 ();
 sky130_fd_sc_hd__decap_3 PHY_10716 ();
 sky130_fd_sc_hd__decap_3 PHY_10717 ();
 sky130_fd_sc_hd__decap_3 PHY_10718 ();
 sky130_fd_sc_hd__decap_3 PHY_10719 ();
 sky130_fd_sc_hd__decap_3 PHY_10720 ();
 sky130_fd_sc_hd__decap_3 PHY_10721 ();
 sky130_fd_sc_hd__decap_3 PHY_10722 ();
 sky130_fd_sc_hd__decap_3 PHY_10723 ();
 sky130_fd_sc_hd__decap_3 PHY_10724 ();
 sky130_fd_sc_hd__decap_3 PHY_10725 ();
 sky130_fd_sc_hd__decap_3 PHY_10726 ();
 sky130_fd_sc_hd__decap_3 PHY_10727 ();
 sky130_fd_sc_hd__decap_3 PHY_10728 ();
 sky130_fd_sc_hd__decap_3 PHY_10729 ();
 sky130_fd_sc_hd__decap_3 PHY_10730 ();
 sky130_fd_sc_hd__decap_3 PHY_10731 ();
 sky130_fd_sc_hd__decap_3 PHY_10732 ();
 sky130_fd_sc_hd__decap_3 PHY_10733 ();
 sky130_fd_sc_hd__decap_3 PHY_10734 ();
 sky130_fd_sc_hd__decap_3 PHY_10735 ();
 sky130_fd_sc_hd__decap_3 PHY_10736 ();
 sky130_fd_sc_hd__decap_3 PHY_10737 ();
 sky130_fd_sc_hd__decap_3 PHY_10738 ();
 sky130_fd_sc_hd__decap_3 PHY_10739 ();
 sky130_fd_sc_hd__decap_3 PHY_10740 ();
 sky130_fd_sc_hd__decap_3 PHY_10741 ();
 sky130_fd_sc_hd__decap_3 PHY_10742 ();
 sky130_fd_sc_hd__decap_3 PHY_10743 ();
 sky130_fd_sc_hd__decap_3 PHY_10744 ();
 sky130_fd_sc_hd__decap_3 PHY_10745 ();
 sky130_fd_sc_hd__decap_3 PHY_10746 ();
 sky130_fd_sc_hd__decap_3 PHY_10747 ();
 sky130_fd_sc_hd__decap_3 PHY_10748 ();
 sky130_fd_sc_hd__decap_3 PHY_10749 ();
 sky130_fd_sc_hd__decap_3 PHY_10750 ();
 sky130_fd_sc_hd__decap_3 PHY_10751 ();
 sky130_fd_sc_hd__decap_3 PHY_10752 ();
 sky130_fd_sc_hd__decap_3 PHY_10753 ();
 sky130_fd_sc_hd__decap_3 PHY_10754 ();
 sky130_fd_sc_hd__decap_3 PHY_10755 ();
 sky130_fd_sc_hd__decap_3 PHY_10756 ();
 sky130_fd_sc_hd__decap_3 PHY_10757 ();
 sky130_fd_sc_hd__decap_3 PHY_10758 ();
 sky130_fd_sc_hd__decap_3 PHY_10759 ();
 sky130_fd_sc_hd__decap_3 PHY_10760 ();
 sky130_fd_sc_hd__decap_3 PHY_10761 ();
 sky130_fd_sc_hd__decap_3 PHY_10762 ();
 sky130_fd_sc_hd__decap_3 PHY_10763 ();
 sky130_fd_sc_hd__decap_3 PHY_10764 ();
 sky130_fd_sc_hd__decap_3 PHY_10765 ();
 sky130_fd_sc_hd__decap_3 PHY_10766 ();
 sky130_fd_sc_hd__decap_3 PHY_10767 ();
 sky130_fd_sc_hd__decap_3 PHY_10768 ();
 sky130_fd_sc_hd__decap_3 PHY_10769 ();
 sky130_fd_sc_hd__decap_3 PHY_10770 ();
 sky130_fd_sc_hd__decap_3 PHY_10771 ();
 sky130_fd_sc_hd__decap_3 PHY_10772 ();
 sky130_fd_sc_hd__decap_3 PHY_10773 ();
 sky130_fd_sc_hd__decap_3 PHY_10774 ();
 sky130_fd_sc_hd__decap_3 PHY_10775 ();
 sky130_fd_sc_hd__decap_3 PHY_10776 ();
 sky130_fd_sc_hd__decap_3 PHY_10777 ();
 sky130_fd_sc_hd__decap_3 PHY_10778 ();
 sky130_fd_sc_hd__decap_3 PHY_10779 ();
 sky130_fd_sc_hd__decap_3 PHY_10780 ();
 sky130_fd_sc_hd__decap_3 PHY_10781 ();
 sky130_fd_sc_hd__decap_3 PHY_10782 ();
 sky130_fd_sc_hd__decap_3 PHY_10783 ();
 sky130_fd_sc_hd__decap_3 PHY_10784 ();
 sky130_fd_sc_hd__decap_3 PHY_10785 ();
 sky130_fd_sc_hd__decap_3 PHY_10786 ();
 sky130_fd_sc_hd__decap_3 PHY_10787 ();
 sky130_fd_sc_hd__decap_3 PHY_10788 ();
 sky130_fd_sc_hd__decap_3 PHY_10789 ();
 sky130_fd_sc_hd__decap_3 PHY_10790 ();
 sky130_fd_sc_hd__decap_3 PHY_10791 ();
 sky130_fd_sc_hd__decap_3 PHY_10792 ();
 sky130_fd_sc_hd__decap_3 PHY_10793 ();
 sky130_fd_sc_hd__decap_3 PHY_10794 ();
 sky130_fd_sc_hd__decap_3 PHY_10795 ();
 sky130_fd_sc_hd__decap_3 PHY_10796 ();
 sky130_fd_sc_hd__decap_3 PHY_10797 ();
 sky130_fd_sc_hd__decap_3 PHY_10798 ();
 sky130_fd_sc_hd__decap_3 PHY_10799 ();
 sky130_fd_sc_hd__decap_3 PHY_10800 ();
 sky130_fd_sc_hd__decap_3 PHY_10801 ();
 sky130_fd_sc_hd__decap_3 PHY_10802 ();
 sky130_fd_sc_hd__decap_3 PHY_10803 ();
 sky130_fd_sc_hd__decap_3 PHY_10804 ();
 sky130_fd_sc_hd__decap_3 PHY_10805 ();
 sky130_fd_sc_hd__decap_3 PHY_10806 ();
 sky130_fd_sc_hd__decap_3 PHY_10807 ();
 sky130_fd_sc_hd__decap_3 PHY_10808 ();
 sky130_fd_sc_hd__decap_3 PHY_10809 ();
 sky130_fd_sc_hd__decap_3 PHY_10810 ();
 sky130_fd_sc_hd__decap_3 PHY_10811 ();
 sky130_fd_sc_hd__decap_3 PHY_10812 ();
 sky130_fd_sc_hd__decap_3 PHY_10813 ();
 sky130_fd_sc_hd__decap_3 PHY_10814 ();
 sky130_fd_sc_hd__decap_3 PHY_10815 ();
 sky130_fd_sc_hd__decap_3 PHY_10816 ();
 sky130_fd_sc_hd__decap_3 PHY_10817 ();
 sky130_fd_sc_hd__decap_3 PHY_10818 ();
 sky130_fd_sc_hd__decap_3 PHY_10819 ();
 sky130_fd_sc_hd__decap_3 PHY_10820 ();
 sky130_fd_sc_hd__decap_3 PHY_10821 ();
 sky130_fd_sc_hd__decap_3 PHY_10822 ();
 sky130_fd_sc_hd__decap_3 PHY_10823 ();
 sky130_fd_sc_hd__decap_3 PHY_10824 ();
 sky130_fd_sc_hd__decap_3 PHY_10825 ();
 sky130_fd_sc_hd__decap_3 PHY_10826 ();
 sky130_fd_sc_hd__decap_3 PHY_10827 ();
 sky130_fd_sc_hd__decap_3 PHY_10828 ();
 sky130_fd_sc_hd__decap_3 PHY_10829 ();
 sky130_fd_sc_hd__decap_3 PHY_10830 ();
 sky130_fd_sc_hd__decap_3 PHY_10831 ();
 sky130_fd_sc_hd__decap_3 PHY_10832 ();
 sky130_fd_sc_hd__decap_3 PHY_10833 ();
 sky130_fd_sc_hd__decap_3 PHY_10834 ();
 sky130_fd_sc_hd__decap_3 PHY_10835 ();
 sky130_fd_sc_hd__decap_3 PHY_10836 ();
 sky130_fd_sc_hd__decap_3 PHY_10837 ();
 sky130_fd_sc_hd__decap_3 PHY_10838 ();
 sky130_fd_sc_hd__decap_3 PHY_10839 ();
 sky130_fd_sc_hd__decap_3 PHY_10840 ();
 sky130_fd_sc_hd__decap_3 PHY_10841 ();
 sky130_fd_sc_hd__decap_3 PHY_10842 ();
 sky130_fd_sc_hd__decap_3 PHY_10843 ();
 sky130_fd_sc_hd__decap_3 PHY_10844 ();
 sky130_fd_sc_hd__decap_3 PHY_10845 ();
 sky130_fd_sc_hd__decap_3 PHY_10846 ();
 sky130_fd_sc_hd__decap_3 PHY_10847 ();
 sky130_fd_sc_hd__decap_3 PHY_10848 ();
 sky130_fd_sc_hd__decap_3 PHY_10849 ();
 sky130_fd_sc_hd__decap_3 PHY_10850 ();
 sky130_fd_sc_hd__decap_3 PHY_10851 ();
 sky130_fd_sc_hd__decap_3 PHY_10852 ();
 sky130_fd_sc_hd__decap_3 PHY_10853 ();
 sky130_fd_sc_hd__decap_3 PHY_10854 ();
 sky130_fd_sc_hd__decap_3 PHY_10855 ();
 sky130_fd_sc_hd__decap_3 PHY_10856 ();
 sky130_fd_sc_hd__decap_3 PHY_10857 ();
 sky130_fd_sc_hd__decap_3 PHY_10858 ();
 sky130_fd_sc_hd__decap_3 PHY_10859 ();
 sky130_fd_sc_hd__decap_3 PHY_10860 ();
 sky130_fd_sc_hd__decap_3 PHY_10861 ();
 sky130_fd_sc_hd__decap_3 PHY_10862 ();
 sky130_fd_sc_hd__decap_3 PHY_10863 ();
 sky130_fd_sc_hd__decap_3 PHY_10864 ();
 sky130_fd_sc_hd__decap_3 PHY_10865 ();
 sky130_fd_sc_hd__decap_3 PHY_10866 ();
 sky130_fd_sc_hd__decap_3 PHY_10867 ();
 sky130_fd_sc_hd__decap_3 PHY_10868 ();
 sky130_fd_sc_hd__decap_3 PHY_10869 ();
 sky130_fd_sc_hd__decap_3 PHY_10870 ();
 sky130_fd_sc_hd__decap_3 PHY_10871 ();
 sky130_fd_sc_hd__decap_3 PHY_10872 ();
 sky130_fd_sc_hd__decap_3 PHY_10873 ();
 sky130_fd_sc_hd__decap_3 PHY_10874 ();
 sky130_fd_sc_hd__decap_3 PHY_10875 ();
 sky130_fd_sc_hd__decap_3 PHY_10876 ();
 sky130_fd_sc_hd__decap_3 PHY_10877 ();
 sky130_fd_sc_hd__decap_3 PHY_10878 ();
 sky130_fd_sc_hd__decap_3 PHY_10879 ();
 sky130_fd_sc_hd__decap_3 PHY_10880 ();
 sky130_fd_sc_hd__decap_3 PHY_10881 ();
 sky130_fd_sc_hd__decap_3 PHY_10882 ();
 sky130_fd_sc_hd__decap_3 PHY_10883 ();
 sky130_fd_sc_hd__decap_3 PHY_10884 ();
 sky130_fd_sc_hd__decap_3 PHY_10885 ();
 sky130_fd_sc_hd__decap_3 PHY_10886 ();
 sky130_fd_sc_hd__decap_3 PHY_10887 ();
 sky130_fd_sc_hd__decap_3 PHY_10888 ();
 sky130_fd_sc_hd__decap_3 PHY_10889 ();
 sky130_fd_sc_hd__decap_3 PHY_10890 ();
 sky130_fd_sc_hd__decap_3 PHY_10891 ();
 sky130_fd_sc_hd__decap_3 PHY_10892 ();
 sky130_fd_sc_hd__decap_3 PHY_10893 ();
 sky130_fd_sc_hd__decap_3 PHY_10894 ();
 sky130_fd_sc_hd__decap_3 PHY_10895 ();
 sky130_fd_sc_hd__decap_3 PHY_10896 ();
 sky130_fd_sc_hd__decap_3 PHY_10897 ();
 sky130_fd_sc_hd__decap_3 PHY_10898 ();
 sky130_fd_sc_hd__decap_3 PHY_10899 ();
 sky130_fd_sc_hd__decap_3 PHY_10900 ();
 sky130_fd_sc_hd__decap_3 PHY_10901 ();
 sky130_fd_sc_hd__decap_3 PHY_10902 ();
 sky130_fd_sc_hd__decap_3 PHY_10903 ();
 sky130_fd_sc_hd__decap_3 PHY_10904 ();
 sky130_fd_sc_hd__decap_3 PHY_10905 ();
 sky130_fd_sc_hd__decap_3 PHY_10906 ();
 sky130_fd_sc_hd__decap_3 PHY_10907 ();
 sky130_fd_sc_hd__decap_3 PHY_10908 ();
 sky130_fd_sc_hd__decap_3 PHY_10909 ();
 sky130_fd_sc_hd__decap_3 PHY_10910 ();
 sky130_fd_sc_hd__decap_3 PHY_10911 ();
 sky130_fd_sc_hd__decap_3 PHY_10912 ();
 sky130_fd_sc_hd__decap_3 PHY_10913 ();
 sky130_fd_sc_hd__decap_3 PHY_10914 ();
 sky130_fd_sc_hd__decap_3 PHY_10915 ();
 sky130_fd_sc_hd__decap_3 PHY_10916 ();
 sky130_fd_sc_hd__decap_3 PHY_10917 ();
 sky130_fd_sc_hd__decap_3 PHY_10918 ();
 sky130_fd_sc_hd__decap_3 PHY_10919 ();
 sky130_fd_sc_hd__decap_3 PHY_10920 ();
 sky130_fd_sc_hd__decap_3 PHY_10921 ();
 sky130_fd_sc_hd__decap_3 PHY_10922 ();
 sky130_fd_sc_hd__decap_3 PHY_10923 ();
 sky130_fd_sc_hd__decap_3 PHY_10924 ();
 sky130_fd_sc_hd__decap_3 PHY_10925 ();
 sky130_fd_sc_hd__decap_3 PHY_10926 ();
 sky130_fd_sc_hd__decap_3 PHY_10927 ();
 sky130_fd_sc_hd__decap_3 PHY_10928 ();
 sky130_fd_sc_hd__decap_3 PHY_10929 ();
 sky130_fd_sc_hd__decap_3 PHY_10930 ();
 sky130_fd_sc_hd__decap_3 PHY_10931 ();
 sky130_fd_sc_hd__decap_3 PHY_10932 ();
 sky130_fd_sc_hd__decap_3 PHY_10933 ();
 sky130_fd_sc_hd__decap_3 PHY_10934 ();
 sky130_fd_sc_hd__decap_3 PHY_10935 ();
 sky130_fd_sc_hd__decap_3 PHY_10936 ();
 sky130_fd_sc_hd__decap_3 PHY_10937 ();
 sky130_fd_sc_hd__decap_3 PHY_10938 ();
 sky130_fd_sc_hd__decap_3 PHY_10939 ();
 sky130_fd_sc_hd__decap_3 PHY_10940 ();
 sky130_fd_sc_hd__decap_3 PHY_10941 ();
 sky130_fd_sc_hd__decap_3 PHY_10942 ();
 sky130_fd_sc_hd__decap_3 PHY_10943 ();
 sky130_fd_sc_hd__decap_3 PHY_10944 ();
 sky130_fd_sc_hd__decap_3 PHY_10945 ();
 sky130_fd_sc_hd__decap_3 PHY_10946 ();
 sky130_fd_sc_hd__decap_3 PHY_10947 ();
 sky130_fd_sc_hd__decap_3 PHY_10948 ();
 sky130_fd_sc_hd__decap_3 PHY_10949 ();
 sky130_fd_sc_hd__decap_3 PHY_10950 ();
 sky130_fd_sc_hd__decap_3 PHY_10951 ();
 sky130_fd_sc_hd__decap_3 PHY_10952 ();
 sky130_fd_sc_hd__decap_3 PHY_10953 ();
 sky130_fd_sc_hd__decap_3 PHY_10954 ();
 sky130_fd_sc_hd__decap_3 PHY_10955 ();
 sky130_fd_sc_hd__decap_3 PHY_10956 ();
 sky130_fd_sc_hd__decap_3 PHY_10957 ();
 sky130_fd_sc_hd__decap_3 PHY_10958 ();
 sky130_fd_sc_hd__decap_3 PHY_10959 ();
 sky130_fd_sc_hd__decap_3 PHY_10960 ();
 sky130_fd_sc_hd__decap_3 PHY_10961 ();
 sky130_fd_sc_hd__decap_3 PHY_10962 ();
 sky130_fd_sc_hd__decap_3 PHY_10963 ();
 sky130_fd_sc_hd__decap_3 PHY_10964 ();
 sky130_fd_sc_hd__decap_3 PHY_10965 ();
 sky130_fd_sc_hd__decap_3 PHY_10966 ();
 sky130_fd_sc_hd__decap_3 PHY_10967 ();
 sky130_fd_sc_hd__decap_3 PHY_10968 ();
 sky130_fd_sc_hd__decap_3 PHY_10969 ();
 sky130_fd_sc_hd__decap_3 PHY_10970 ();
 sky130_fd_sc_hd__decap_3 PHY_10971 ();
 sky130_fd_sc_hd__decap_3 PHY_10972 ();
 sky130_fd_sc_hd__decap_3 PHY_10973 ();
 sky130_fd_sc_hd__decap_3 PHY_10974 ();
 sky130_fd_sc_hd__decap_3 PHY_10975 ();
 sky130_fd_sc_hd__decap_3 PHY_10976 ();
 sky130_fd_sc_hd__decap_3 PHY_10977 ();
 sky130_fd_sc_hd__decap_3 PHY_10978 ();
 sky130_fd_sc_hd__decap_3 PHY_10979 ();
 sky130_fd_sc_hd__decap_3 PHY_10980 ();
 sky130_fd_sc_hd__decap_3 PHY_10981 ();
 sky130_fd_sc_hd__decap_3 PHY_10982 ();
 sky130_fd_sc_hd__decap_3 PHY_10983 ();
 sky130_fd_sc_hd__decap_3 PHY_10984 ();
 sky130_fd_sc_hd__decap_3 PHY_10985 ();
 sky130_fd_sc_hd__decap_3 PHY_10986 ();
 sky130_fd_sc_hd__decap_3 PHY_10987 ();
 sky130_fd_sc_hd__decap_3 PHY_10988 ();
 sky130_fd_sc_hd__decap_3 PHY_10989 ();
 sky130_fd_sc_hd__decap_3 PHY_10990 ();
 sky130_fd_sc_hd__decap_3 PHY_10991 ();
 sky130_fd_sc_hd__decap_3 PHY_10992 ();
 sky130_fd_sc_hd__decap_3 PHY_10993 ();
 sky130_fd_sc_hd__decap_3 PHY_10994 ();
 sky130_fd_sc_hd__decap_3 PHY_10995 ();
 sky130_fd_sc_hd__decap_3 PHY_10996 ();
 sky130_fd_sc_hd__decap_3 PHY_10997 ();
 sky130_fd_sc_hd__decap_3 PHY_10998 ();
 sky130_fd_sc_hd__decap_3 PHY_10999 ();
 sky130_fd_sc_hd__decap_3 PHY_11000 ();
 sky130_fd_sc_hd__decap_3 PHY_11001 ();
 sky130_fd_sc_hd__decap_3 PHY_11002 ();
 sky130_fd_sc_hd__decap_3 PHY_11003 ();
 sky130_fd_sc_hd__decap_3 PHY_11004 ();
 sky130_fd_sc_hd__decap_3 PHY_11005 ();
 sky130_fd_sc_hd__decap_3 PHY_11006 ();
 sky130_fd_sc_hd__decap_3 PHY_11007 ();
 sky130_fd_sc_hd__decap_3 PHY_11008 ();
 sky130_fd_sc_hd__decap_3 PHY_11009 ();
 sky130_fd_sc_hd__decap_3 PHY_11010 ();
 sky130_fd_sc_hd__decap_3 PHY_11011 ();
 sky130_fd_sc_hd__decap_3 PHY_11012 ();
 sky130_fd_sc_hd__decap_3 PHY_11013 ();
 sky130_fd_sc_hd__decap_3 PHY_11014 ();
 sky130_fd_sc_hd__decap_3 PHY_11015 ();
 sky130_fd_sc_hd__decap_3 PHY_11016 ();
 sky130_fd_sc_hd__decap_3 PHY_11017 ();
 sky130_fd_sc_hd__decap_3 PHY_11018 ();
 sky130_fd_sc_hd__decap_3 PHY_11019 ();
 sky130_fd_sc_hd__decap_3 PHY_11020 ();
 sky130_fd_sc_hd__decap_3 PHY_11021 ();
 sky130_fd_sc_hd__decap_3 PHY_11022 ();
 sky130_fd_sc_hd__decap_3 PHY_11023 ();
 sky130_fd_sc_hd__decap_3 PHY_11024 ();
 sky130_fd_sc_hd__decap_3 PHY_11025 ();
 sky130_fd_sc_hd__decap_3 PHY_11026 ();
 sky130_fd_sc_hd__decap_3 PHY_11027 ();
 sky130_fd_sc_hd__decap_3 PHY_11028 ();
 sky130_fd_sc_hd__decap_3 PHY_11029 ();
 sky130_fd_sc_hd__decap_3 PHY_11030 ();
 sky130_fd_sc_hd__decap_3 PHY_11031 ();
 sky130_fd_sc_hd__decap_3 PHY_11032 ();
 sky130_fd_sc_hd__decap_3 PHY_11033 ();
 sky130_fd_sc_hd__decap_3 PHY_11034 ();
 sky130_fd_sc_hd__decap_3 PHY_11035 ();
 sky130_fd_sc_hd__decap_3 PHY_11036 ();
 sky130_fd_sc_hd__decap_3 PHY_11037 ();
 sky130_fd_sc_hd__decap_3 PHY_11038 ();
 sky130_fd_sc_hd__decap_3 PHY_11039 ();
 sky130_fd_sc_hd__decap_3 PHY_11040 ();
 sky130_fd_sc_hd__decap_3 PHY_11041 ();
 sky130_fd_sc_hd__decap_3 PHY_11042 ();
 sky130_fd_sc_hd__decap_3 PHY_11043 ();
 sky130_fd_sc_hd__decap_3 PHY_11044 ();
 sky130_fd_sc_hd__decap_3 PHY_11045 ();
 sky130_fd_sc_hd__decap_3 PHY_11046 ();
 sky130_fd_sc_hd__decap_3 PHY_11047 ();
 sky130_fd_sc_hd__decap_3 PHY_11048 ();
 sky130_fd_sc_hd__decap_3 PHY_11049 ();
 sky130_fd_sc_hd__decap_3 PHY_11050 ();
 sky130_fd_sc_hd__decap_3 PHY_11051 ();
 sky130_fd_sc_hd__decap_3 PHY_11052 ();
 sky130_fd_sc_hd__decap_3 PHY_11053 ();
 sky130_fd_sc_hd__decap_3 PHY_11054 ();
 sky130_fd_sc_hd__decap_3 PHY_11055 ();
 sky130_fd_sc_hd__decap_3 PHY_11056 ();
 sky130_fd_sc_hd__decap_3 PHY_11057 ();
 sky130_fd_sc_hd__decap_3 PHY_11058 ();
 sky130_fd_sc_hd__decap_3 PHY_11059 ();
 sky130_fd_sc_hd__decap_3 PHY_11060 ();
 sky130_fd_sc_hd__decap_3 PHY_11061 ();
 sky130_fd_sc_hd__decap_3 PHY_11062 ();
 sky130_fd_sc_hd__decap_3 PHY_11063 ();
 sky130_fd_sc_hd__decap_3 PHY_11064 ();
 sky130_fd_sc_hd__decap_3 PHY_11065 ();
 sky130_fd_sc_hd__decap_3 PHY_11066 ();
 sky130_fd_sc_hd__decap_3 PHY_11067 ();
 sky130_fd_sc_hd__decap_3 PHY_11068 ();
 sky130_fd_sc_hd__decap_3 PHY_11069 ();
 sky130_fd_sc_hd__decap_3 PHY_11070 ();
 sky130_fd_sc_hd__decap_3 PHY_11071 ();
 sky130_fd_sc_hd__decap_3 PHY_11072 ();
 sky130_fd_sc_hd__decap_3 PHY_11073 ();
 sky130_fd_sc_hd__decap_3 PHY_11074 ();
 sky130_fd_sc_hd__decap_3 PHY_11075 ();
 sky130_fd_sc_hd__decap_3 PHY_11076 ();
 sky130_fd_sc_hd__decap_3 PHY_11077 ();
 sky130_fd_sc_hd__decap_3 PHY_11078 ();
 sky130_fd_sc_hd__decap_3 PHY_11079 ();
 sky130_fd_sc_hd__decap_3 PHY_11080 ();
 sky130_fd_sc_hd__decap_3 PHY_11081 ();
 sky130_fd_sc_hd__decap_3 PHY_11082 ();
 sky130_fd_sc_hd__decap_3 PHY_11083 ();
 sky130_fd_sc_hd__decap_3 PHY_11084 ();
 sky130_fd_sc_hd__decap_3 PHY_11085 ();
 sky130_fd_sc_hd__decap_3 PHY_11086 ();
 sky130_fd_sc_hd__decap_3 PHY_11087 ();
 sky130_fd_sc_hd__decap_3 PHY_11088 ();
 sky130_fd_sc_hd__decap_3 PHY_11089 ();
 sky130_fd_sc_hd__decap_3 PHY_11090 ();
 sky130_fd_sc_hd__decap_3 PHY_11091 ();
 sky130_fd_sc_hd__decap_3 PHY_11092 ();
 sky130_fd_sc_hd__decap_3 PHY_11093 ();
 sky130_fd_sc_hd__decap_3 PHY_11094 ();
 sky130_fd_sc_hd__decap_3 PHY_11095 ();
 sky130_fd_sc_hd__decap_3 PHY_11096 ();
 sky130_fd_sc_hd__decap_3 PHY_11097 ();
 sky130_fd_sc_hd__decap_3 PHY_11098 ();
 sky130_fd_sc_hd__decap_3 PHY_11099 ();
 sky130_fd_sc_hd__decap_3 PHY_11100 ();
 sky130_fd_sc_hd__decap_3 PHY_11101 ();
 sky130_fd_sc_hd__decap_3 PHY_11102 ();
 sky130_fd_sc_hd__decap_3 PHY_11103 ();
 sky130_fd_sc_hd__decap_3 PHY_11104 ();
 sky130_fd_sc_hd__decap_3 PHY_11105 ();
 sky130_fd_sc_hd__decap_3 PHY_11106 ();
 sky130_fd_sc_hd__decap_3 PHY_11107 ();
 sky130_fd_sc_hd__decap_3 PHY_11108 ();
 sky130_fd_sc_hd__decap_3 PHY_11109 ();
 sky130_fd_sc_hd__decap_3 PHY_11110 ();
 sky130_fd_sc_hd__decap_3 PHY_11111 ();
 sky130_fd_sc_hd__decap_3 PHY_11112 ();
 sky130_fd_sc_hd__decap_3 PHY_11113 ();
 sky130_fd_sc_hd__decap_3 PHY_11114 ();
 sky130_fd_sc_hd__decap_3 PHY_11115 ();
 sky130_fd_sc_hd__decap_3 PHY_11116 ();
 sky130_fd_sc_hd__decap_3 PHY_11117 ();
 sky130_fd_sc_hd__decap_3 PHY_11118 ();
 sky130_fd_sc_hd__decap_3 PHY_11119 ();
 sky130_fd_sc_hd__decap_3 PHY_11120 ();
 sky130_fd_sc_hd__decap_3 PHY_11121 ();
 sky130_fd_sc_hd__decap_3 PHY_11122 ();
 sky130_fd_sc_hd__decap_3 PHY_11123 ();
 sky130_fd_sc_hd__decap_3 PHY_11124 ();
 sky130_fd_sc_hd__decap_3 PHY_11125 ();
 sky130_fd_sc_hd__decap_3 PHY_11126 ();
 sky130_fd_sc_hd__decap_3 PHY_11127 ();
 sky130_fd_sc_hd__decap_3 PHY_11128 ();
 sky130_fd_sc_hd__decap_3 PHY_11129 ();
 sky130_fd_sc_hd__decap_3 PHY_11130 ();
 sky130_fd_sc_hd__decap_3 PHY_11131 ();
 sky130_fd_sc_hd__decap_3 PHY_11132 ();
 sky130_fd_sc_hd__decap_3 PHY_11133 ();
 sky130_fd_sc_hd__decap_3 PHY_11134 ();
 sky130_fd_sc_hd__decap_3 PHY_11135 ();
 sky130_fd_sc_hd__decap_3 PHY_11136 ();
 sky130_fd_sc_hd__decap_3 PHY_11137 ();
 sky130_fd_sc_hd__decap_3 PHY_11138 ();
 sky130_fd_sc_hd__decap_3 PHY_11139 ();
 sky130_fd_sc_hd__decap_3 PHY_11140 ();
 sky130_fd_sc_hd__decap_3 PHY_11141 ();
 sky130_fd_sc_hd__decap_3 PHY_11142 ();
 sky130_fd_sc_hd__decap_3 PHY_11143 ();
 sky130_fd_sc_hd__decap_3 PHY_11144 ();
 sky130_fd_sc_hd__decap_3 PHY_11145 ();
 sky130_fd_sc_hd__decap_3 PHY_11146 ();
 sky130_fd_sc_hd__decap_3 PHY_11147 ();
 sky130_fd_sc_hd__decap_3 PHY_11148 ();
 sky130_fd_sc_hd__decap_3 PHY_11149 ();
 sky130_fd_sc_hd__decap_3 PHY_11150 ();
 sky130_fd_sc_hd__decap_3 PHY_11151 ();
 sky130_fd_sc_hd__decap_3 PHY_11152 ();
 sky130_fd_sc_hd__decap_3 PHY_11153 ();
 sky130_fd_sc_hd__decap_3 PHY_11154 ();
 sky130_fd_sc_hd__decap_3 PHY_11155 ();
 sky130_fd_sc_hd__decap_3 PHY_11156 ();
 sky130_fd_sc_hd__decap_3 PHY_11157 ();
 sky130_fd_sc_hd__decap_3 PHY_11158 ();
 sky130_fd_sc_hd__decap_3 PHY_11159 ();
 sky130_fd_sc_hd__decap_3 PHY_11160 ();
 sky130_fd_sc_hd__decap_3 PHY_11161 ();
 sky130_fd_sc_hd__decap_3 PHY_11162 ();
 sky130_fd_sc_hd__decap_3 PHY_11163 ();
 sky130_fd_sc_hd__decap_3 PHY_11164 ();
 sky130_fd_sc_hd__decap_3 PHY_11165 ();
 sky130_fd_sc_hd__decap_3 PHY_11166 ();
 sky130_fd_sc_hd__decap_3 PHY_11167 ();
 sky130_fd_sc_hd__decap_3 PHY_11168 ();
 sky130_fd_sc_hd__decap_3 PHY_11169 ();
 sky130_fd_sc_hd__decap_3 PHY_11170 ();
 sky130_fd_sc_hd__decap_3 PHY_11171 ();
 sky130_fd_sc_hd__decap_3 PHY_11172 ();
 sky130_fd_sc_hd__decap_3 PHY_11173 ();
 sky130_fd_sc_hd__decap_3 PHY_11174 ();
 sky130_fd_sc_hd__decap_3 PHY_11175 ();
 sky130_fd_sc_hd__decap_3 PHY_11176 ();
 sky130_fd_sc_hd__decap_3 PHY_11177 ();
 sky130_fd_sc_hd__decap_3 PHY_11178 ();
 sky130_fd_sc_hd__decap_3 PHY_11179 ();
 sky130_fd_sc_hd__decap_3 PHY_11180 ();
 sky130_fd_sc_hd__decap_3 PHY_11181 ();
 sky130_fd_sc_hd__decap_3 PHY_11182 ();
 sky130_fd_sc_hd__decap_3 PHY_11183 ();
 sky130_fd_sc_hd__decap_3 PHY_11184 ();
 sky130_fd_sc_hd__decap_3 PHY_11185 ();
 sky130_fd_sc_hd__decap_3 PHY_11186 ();
 sky130_fd_sc_hd__decap_3 PHY_11187 ();
 sky130_fd_sc_hd__decap_3 PHY_11188 ();
 sky130_fd_sc_hd__decap_3 PHY_11189 ();
 sky130_fd_sc_hd__decap_3 PHY_11190 ();
 sky130_fd_sc_hd__decap_3 PHY_11191 ();
 sky130_fd_sc_hd__decap_3 PHY_11192 ();
 sky130_fd_sc_hd__decap_3 PHY_11193 ();
 sky130_fd_sc_hd__decap_3 PHY_11194 ();
 sky130_fd_sc_hd__decap_3 PHY_11195 ();
 sky130_fd_sc_hd__decap_3 PHY_11196 ();
 sky130_fd_sc_hd__decap_3 PHY_11197 ();
 sky130_fd_sc_hd__decap_3 PHY_11198 ();
 sky130_fd_sc_hd__decap_3 PHY_11199 ();
 sky130_fd_sc_hd__decap_3 PHY_11200 ();
 sky130_fd_sc_hd__decap_3 PHY_11201 ();
 sky130_fd_sc_hd__decap_3 PHY_11202 ();
 sky130_fd_sc_hd__decap_3 PHY_11203 ();
 sky130_fd_sc_hd__decap_3 PHY_11204 ();
 sky130_fd_sc_hd__decap_3 PHY_11205 ();
 sky130_fd_sc_hd__decap_3 PHY_11206 ();
 sky130_fd_sc_hd__decap_3 PHY_11207 ();
 sky130_fd_sc_hd__decap_3 PHY_11208 ();
 sky130_fd_sc_hd__decap_3 PHY_11209 ();
 sky130_fd_sc_hd__decap_3 PHY_11210 ();
 sky130_fd_sc_hd__decap_3 PHY_11211 ();
 sky130_fd_sc_hd__decap_3 PHY_11212 ();
 sky130_fd_sc_hd__decap_3 PHY_11213 ();
 sky130_fd_sc_hd__decap_3 PHY_11214 ();
 sky130_fd_sc_hd__decap_3 PHY_11215 ();
 sky130_fd_sc_hd__decap_3 PHY_11216 ();
 sky130_fd_sc_hd__decap_3 PHY_11217 ();
 sky130_fd_sc_hd__decap_3 PHY_11218 ();
 sky130_fd_sc_hd__decap_3 PHY_11219 ();
 sky130_fd_sc_hd__decap_3 PHY_11220 ();
 sky130_fd_sc_hd__decap_3 PHY_11221 ();
 sky130_fd_sc_hd__decap_3 PHY_11222 ();
 sky130_fd_sc_hd__decap_3 PHY_11223 ();
 sky130_fd_sc_hd__decap_3 PHY_11224 ();
 sky130_fd_sc_hd__decap_3 PHY_11225 ();
 sky130_fd_sc_hd__decap_3 PHY_11226 ();
 sky130_fd_sc_hd__decap_3 PHY_11227 ();
 sky130_fd_sc_hd__decap_3 PHY_11228 ();
 sky130_fd_sc_hd__decap_3 PHY_11229 ();
 sky130_fd_sc_hd__decap_3 PHY_11230 ();
 sky130_fd_sc_hd__decap_3 PHY_11231 ();
 sky130_fd_sc_hd__decap_3 PHY_11232 ();
 sky130_fd_sc_hd__decap_3 PHY_11233 ();
 sky130_fd_sc_hd__decap_3 PHY_11234 ();
 sky130_fd_sc_hd__decap_3 PHY_11235 ();
 sky130_fd_sc_hd__decap_3 PHY_11236 ();
 sky130_fd_sc_hd__decap_3 PHY_11237 ();
 sky130_fd_sc_hd__decap_3 PHY_11238 ();
 sky130_fd_sc_hd__decap_3 PHY_11239 ();
 sky130_fd_sc_hd__decap_3 PHY_11240 ();
 sky130_fd_sc_hd__decap_3 PHY_11241 ();
 sky130_fd_sc_hd__decap_3 PHY_11242 ();
 sky130_fd_sc_hd__decap_3 PHY_11243 ();
 sky130_fd_sc_hd__decap_3 PHY_11244 ();
 sky130_fd_sc_hd__decap_3 PHY_11245 ();
 sky130_fd_sc_hd__decap_3 PHY_11246 ();
 sky130_fd_sc_hd__decap_3 PHY_11247 ();
 sky130_fd_sc_hd__decap_3 PHY_11248 ();
 sky130_fd_sc_hd__decap_3 PHY_11249 ();
 sky130_fd_sc_hd__decap_3 PHY_11250 ();
 sky130_fd_sc_hd__decap_3 PHY_11251 ();
 sky130_fd_sc_hd__decap_3 PHY_11252 ();
 sky130_fd_sc_hd__decap_3 PHY_11253 ();
 sky130_fd_sc_hd__decap_3 PHY_11254 ();
 sky130_fd_sc_hd__decap_3 PHY_11255 ();
 sky130_fd_sc_hd__decap_3 PHY_11256 ();
 sky130_fd_sc_hd__decap_3 PHY_11257 ();
 sky130_fd_sc_hd__decap_3 PHY_11258 ();
 sky130_fd_sc_hd__decap_3 PHY_11259 ();
 sky130_fd_sc_hd__decap_3 PHY_11260 ();
 sky130_fd_sc_hd__decap_3 PHY_11261 ();
 sky130_fd_sc_hd__decap_3 PHY_11262 ();
 sky130_fd_sc_hd__decap_3 PHY_11263 ();
 sky130_fd_sc_hd__decap_3 PHY_11264 ();
 sky130_fd_sc_hd__decap_3 PHY_11265 ();
 sky130_fd_sc_hd__decap_3 PHY_11266 ();
 sky130_fd_sc_hd__decap_3 PHY_11267 ();
 sky130_fd_sc_hd__decap_3 PHY_11268 ();
 sky130_fd_sc_hd__decap_3 PHY_11269 ();
 sky130_fd_sc_hd__decap_3 PHY_11270 ();
 sky130_fd_sc_hd__decap_3 PHY_11271 ();
 sky130_fd_sc_hd__decap_3 PHY_11272 ();
 sky130_fd_sc_hd__decap_3 PHY_11273 ();
 sky130_fd_sc_hd__decap_3 PHY_11274 ();
 sky130_fd_sc_hd__decap_3 PHY_11275 ();
 sky130_fd_sc_hd__decap_3 PHY_11276 ();
 sky130_fd_sc_hd__decap_3 PHY_11277 ();
 sky130_fd_sc_hd__decap_3 PHY_11278 ();
 sky130_fd_sc_hd__decap_3 PHY_11279 ();
 sky130_fd_sc_hd__decap_3 PHY_11280 ();
 sky130_fd_sc_hd__decap_3 PHY_11281 ();
 sky130_fd_sc_hd__decap_3 PHY_11282 ();
 sky130_fd_sc_hd__decap_3 PHY_11283 ();
 sky130_fd_sc_hd__decap_3 PHY_11284 ();
 sky130_fd_sc_hd__decap_3 PHY_11285 ();
 sky130_fd_sc_hd__decap_3 PHY_11286 ();
 sky130_fd_sc_hd__decap_3 PHY_11287 ();
 sky130_fd_sc_hd__decap_3 PHY_11288 ();
 sky130_fd_sc_hd__decap_3 PHY_11289 ();
 sky130_fd_sc_hd__decap_3 PHY_11290 ();
 sky130_fd_sc_hd__decap_3 PHY_11291 ();
 sky130_fd_sc_hd__decap_3 PHY_11292 ();
 sky130_fd_sc_hd__decap_3 PHY_11293 ();
 sky130_fd_sc_hd__decap_3 PHY_11294 ();
 sky130_fd_sc_hd__decap_3 PHY_11295 ();
 sky130_fd_sc_hd__decap_3 PHY_11296 ();
 sky130_fd_sc_hd__decap_3 PHY_11297 ();
 sky130_fd_sc_hd__decap_3 PHY_11298 ();
 sky130_fd_sc_hd__decap_3 PHY_11299 ();
 sky130_fd_sc_hd__decap_3 PHY_11300 ();
 sky130_fd_sc_hd__decap_3 PHY_11301 ();
 sky130_fd_sc_hd__decap_3 PHY_11302 ();
 sky130_fd_sc_hd__decap_3 PHY_11303 ();
 sky130_fd_sc_hd__decap_3 PHY_11304 ();
 sky130_fd_sc_hd__decap_3 PHY_11305 ();
 sky130_fd_sc_hd__decap_3 PHY_11306 ();
 sky130_fd_sc_hd__decap_3 PHY_11307 ();
 sky130_fd_sc_hd__decap_3 PHY_11308 ();
 sky130_fd_sc_hd__decap_3 PHY_11309 ();
 sky130_fd_sc_hd__decap_3 PHY_11310 ();
 sky130_fd_sc_hd__decap_3 PHY_11311 ();
 sky130_fd_sc_hd__decap_3 PHY_11312 ();
 sky130_fd_sc_hd__decap_3 PHY_11313 ();
 sky130_fd_sc_hd__decap_3 PHY_11314 ();
 sky130_fd_sc_hd__decap_3 PHY_11315 ();
 sky130_fd_sc_hd__decap_3 PHY_11316 ();
 sky130_fd_sc_hd__decap_3 PHY_11317 ();
 sky130_fd_sc_hd__decap_3 PHY_11318 ();
 sky130_fd_sc_hd__decap_3 PHY_11319 ();
 sky130_fd_sc_hd__decap_3 PHY_11320 ();
 sky130_fd_sc_hd__decap_3 PHY_11321 ();
 sky130_fd_sc_hd__decap_3 PHY_11322 ();
 sky130_fd_sc_hd__decap_3 PHY_11323 ();
 sky130_fd_sc_hd__decap_3 PHY_11324 ();
 sky130_fd_sc_hd__decap_3 PHY_11325 ();
 sky130_fd_sc_hd__decap_3 PHY_11326 ();
 sky130_fd_sc_hd__decap_3 PHY_11327 ();
 sky130_fd_sc_hd__decap_3 PHY_11328 ();
 sky130_fd_sc_hd__decap_3 PHY_11329 ();
 sky130_fd_sc_hd__decap_3 PHY_11330 ();
 sky130_fd_sc_hd__decap_3 PHY_11331 ();
 sky130_fd_sc_hd__decap_3 PHY_11332 ();
 sky130_fd_sc_hd__decap_3 PHY_11333 ();
 sky130_fd_sc_hd__decap_3 PHY_11334 ();
 sky130_fd_sc_hd__decap_3 PHY_11335 ();
 sky130_fd_sc_hd__decap_3 PHY_11336 ();
 sky130_fd_sc_hd__decap_3 PHY_11337 ();
 sky130_fd_sc_hd__decap_3 PHY_11338 ();
 sky130_fd_sc_hd__decap_3 PHY_11339 ();
 sky130_fd_sc_hd__decap_3 PHY_11340 ();
 sky130_fd_sc_hd__decap_3 PHY_11341 ();
 sky130_fd_sc_hd__decap_3 PHY_11342 ();
 sky130_fd_sc_hd__decap_3 PHY_11343 ();
 sky130_fd_sc_hd__decap_3 PHY_11344 ();
 sky130_fd_sc_hd__decap_3 PHY_11345 ();
 sky130_fd_sc_hd__decap_3 PHY_11346 ();
 sky130_fd_sc_hd__decap_3 PHY_11347 ();
 sky130_fd_sc_hd__decap_3 PHY_11348 ();
 sky130_fd_sc_hd__decap_3 PHY_11349 ();
 sky130_fd_sc_hd__decap_3 PHY_11350 ();
 sky130_fd_sc_hd__decap_3 PHY_11351 ();
 sky130_fd_sc_hd__decap_3 PHY_11352 ();
 sky130_fd_sc_hd__decap_3 PHY_11353 ();
 sky130_fd_sc_hd__decap_3 PHY_11354 ();
 sky130_fd_sc_hd__decap_3 PHY_11355 ();
 sky130_fd_sc_hd__decap_3 PHY_11356 ();
 sky130_fd_sc_hd__decap_3 PHY_11357 ();
 sky130_fd_sc_hd__decap_3 PHY_11358 ();
 sky130_fd_sc_hd__decap_3 PHY_11359 ();
 sky130_fd_sc_hd__decap_3 PHY_11360 ();
 sky130_fd_sc_hd__decap_3 PHY_11361 ();
 sky130_fd_sc_hd__decap_3 PHY_11362 ();
 sky130_fd_sc_hd__decap_3 PHY_11363 ();
 sky130_fd_sc_hd__decap_3 PHY_11364 ();
 sky130_fd_sc_hd__decap_3 PHY_11365 ();
 sky130_fd_sc_hd__decap_3 PHY_11366 ();
 sky130_fd_sc_hd__decap_3 PHY_11367 ();
 sky130_fd_sc_hd__decap_3 PHY_11368 ();
 sky130_fd_sc_hd__decap_3 PHY_11369 ();
 sky130_fd_sc_hd__decap_3 PHY_11370 ();
 sky130_fd_sc_hd__decap_3 PHY_11371 ();
 sky130_fd_sc_hd__decap_3 PHY_11372 ();
 sky130_fd_sc_hd__decap_3 PHY_11373 ();
 sky130_fd_sc_hd__decap_3 PHY_11374 ();
 sky130_fd_sc_hd__decap_3 PHY_11375 ();
 sky130_fd_sc_hd__decap_3 PHY_11376 ();
 sky130_fd_sc_hd__decap_3 PHY_11377 ();
 sky130_fd_sc_hd__decap_3 PHY_11378 ();
 sky130_fd_sc_hd__decap_3 PHY_11379 ();
 sky130_fd_sc_hd__decap_3 PHY_11380 ();
 sky130_fd_sc_hd__decap_3 PHY_11381 ();
 sky130_fd_sc_hd__decap_3 PHY_11382 ();
 sky130_fd_sc_hd__decap_3 PHY_11383 ();
 sky130_fd_sc_hd__decap_3 PHY_11384 ();
 sky130_fd_sc_hd__decap_3 PHY_11385 ();
 sky130_fd_sc_hd__decap_3 PHY_11386 ();
 sky130_fd_sc_hd__decap_3 PHY_11387 ();
 sky130_fd_sc_hd__decap_3 PHY_11388 ();
 sky130_fd_sc_hd__decap_3 PHY_11389 ();
 sky130_fd_sc_hd__decap_3 PHY_11390 ();
 sky130_fd_sc_hd__decap_3 PHY_11391 ();
 sky130_fd_sc_hd__decap_3 PHY_11392 ();
 sky130_fd_sc_hd__decap_3 PHY_11393 ();
 sky130_fd_sc_hd__decap_3 PHY_11394 ();
 sky130_fd_sc_hd__decap_3 PHY_11395 ();
 sky130_fd_sc_hd__decap_3 PHY_11396 ();
 sky130_fd_sc_hd__decap_3 PHY_11397 ();
 sky130_fd_sc_hd__decap_3 PHY_11398 ();
 sky130_fd_sc_hd__decap_3 PHY_11399 ();
 sky130_fd_sc_hd__decap_3 PHY_11400 ();
 sky130_fd_sc_hd__decap_3 PHY_11401 ();
 sky130_fd_sc_hd__decap_3 PHY_11402 ();
 sky130_fd_sc_hd__decap_3 PHY_11403 ();
 sky130_fd_sc_hd__decap_3 PHY_11404 ();
 sky130_fd_sc_hd__decap_3 PHY_11405 ();
 sky130_fd_sc_hd__decap_3 PHY_11406 ();
 sky130_fd_sc_hd__decap_3 PHY_11407 ();
 sky130_fd_sc_hd__decap_3 PHY_11408 ();
 sky130_fd_sc_hd__decap_3 PHY_11409 ();
 sky130_fd_sc_hd__decap_3 PHY_11410 ();
 sky130_fd_sc_hd__decap_3 PHY_11411 ();
 sky130_fd_sc_hd__decap_3 PHY_11412 ();
 sky130_fd_sc_hd__decap_3 PHY_11413 ();
 sky130_fd_sc_hd__decap_3 PHY_11414 ();
 sky130_fd_sc_hd__decap_3 PHY_11415 ();
 sky130_fd_sc_hd__decap_3 PHY_11416 ();
 sky130_fd_sc_hd__decap_3 PHY_11417 ();
 sky130_fd_sc_hd__decap_3 PHY_11418 ();
 sky130_fd_sc_hd__decap_3 PHY_11419 ();
 sky130_fd_sc_hd__decap_3 PHY_11420 ();
 sky130_fd_sc_hd__decap_3 PHY_11421 ();
 sky130_fd_sc_hd__decap_3 PHY_11422 ();
 sky130_fd_sc_hd__decap_3 PHY_11423 ();
 sky130_fd_sc_hd__decap_3 PHY_11424 ();
 sky130_fd_sc_hd__decap_3 PHY_11425 ();
 sky130_fd_sc_hd__decap_3 PHY_11426 ();
 sky130_fd_sc_hd__decap_3 PHY_11427 ();
 sky130_fd_sc_hd__decap_3 PHY_11428 ();
 sky130_fd_sc_hd__decap_3 PHY_11429 ();
 sky130_fd_sc_hd__decap_3 PHY_11430 ();
 sky130_fd_sc_hd__decap_3 PHY_11431 ();
 sky130_fd_sc_hd__decap_3 PHY_11432 ();
 sky130_fd_sc_hd__decap_3 PHY_11433 ();
 sky130_fd_sc_hd__decap_3 PHY_11434 ();
 sky130_fd_sc_hd__decap_3 PHY_11435 ();
 sky130_fd_sc_hd__decap_3 PHY_11436 ();
 sky130_fd_sc_hd__decap_3 PHY_11437 ();
 sky130_fd_sc_hd__decap_3 PHY_11438 ();
 sky130_fd_sc_hd__decap_3 PHY_11439 ();
 sky130_fd_sc_hd__decap_3 PHY_11440 ();
 sky130_fd_sc_hd__decap_3 PHY_11441 ();
 sky130_fd_sc_hd__decap_3 PHY_11442 ();
 sky130_fd_sc_hd__decap_3 PHY_11443 ();
 sky130_fd_sc_hd__decap_3 PHY_11444 ();
 sky130_fd_sc_hd__decap_3 PHY_11445 ();
 sky130_fd_sc_hd__decap_3 PHY_11446 ();
 sky130_fd_sc_hd__decap_3 PHY_11447 ();
 sky130_fd_sc_hd__decap_3 PHY_11448 ();
 sky130_fd_sc_hd__decap_3 PHY_11449 ();
 sky130_fd_sc_hd__decap_3 PHY_11450 ();
 sky130_fd_sc_hd__decap_3 PHY_11451 ();
 sky130_fd_sc_hd__decap_3 PHY_11452 ();
 sky130_fd_sc_hd__decap_3 PHY_11453 ();
 sky130_fd_sc_hd__decap_3 PHY_11454 ();
 sky130_fd_sc_hd__decap_3 PHY_11455 ();
 sky130_fd_sc_hd__decap_3 PHY_11456 ();
 sky130_fd_sc_hd__decap_3 PHY_11457 ();
 sky130_fd_sc_hd__decap_3 PHY_11458 ();
 sky130_fd_sc_hd__decap_3 PHY_11459 ();
 sky130_fd_sc_hd__decap_3 PHY_11460 ();
 sky130_fd_sc_hd__decap_3 PHY_11461 ();
 sky130_fd_sc_hd__decap_3 PHY_11462 ();
 sky130_fd_sc_hd__decap_3 PHY_11463 ();
 sky130_fd_sc_hd__decap_3 PHY_11464 ();
 sky130_fd_sc_hd__decap_3 PHY_11465 ();
 sky130_fd_sc_hd__decap_3 PHY_11466 ();
 sky130_fd_sc_hd__decap_3 PHY_11467 ();
 sky130_fd_sc_hd__decap_3 PHY_11468 ();
 sky130_fd_sc_hd__decap_3 PHY_11469 ();
 sky130_fd_sc_hd__decap_3 PHY_11470 ();
 sky130_fd_sc_hd__decap_3 PHY_11471 ();
 sky130_fd_sc_hd__decap_3 PHY_11472 ();
 sky130_fd_sc_hd__decap_3 PHY_11473 ();
 sky130_fd_sc_hd__decap_3 PHY_11474 ();
 sky130_fd_sc_hd__decap_3 PHY_11475 ();
 sky130_fd_sc_hd__decap_3 PHY_11476 ();
 sky130_fd_sc_hd__decap_3 PHY_11477 ();
 sky130_fd_sc_hd__decap_3 PHY_11478 ();
 sky130_fd_sc_hd__decap_3 PHY_11479 ();
 sky130_fd_sc_hd__decap_3 PHY_11480 ();
 sky130_fd_sc_hd__decap_3 PHY_11481 ();
 sky130_fd_sc_hd__decap_3 PHY_11482 ();
 sky130_fd_sc_hd__decap_3 PHY_11483 ();
 sky130_fd_sc_hd__decap_3 PHY_11484 ();
 sky130_fd_sc_hd__decap_3 PHY_11485 ();
 sky130_fd_sc_hd__decap_3 PHY_11486 ();
 sky130_fd_sc_hd__decap_3 PHY_11487 ();
 sky130_fd_sc_hd__decap_3 PHY_11488 ();
 sky130_fd_sc_hd__decap_3 PHY_11489 ();
 sky130_fd_sc_hd__decap_3 PHY_11490 ();
 sky130_fd_sc_hd__decap_3 PHY_11491 ();
 sky130_fd_sc_hd__decap_3 PHY_11492 ();
 sky130_fd_sc_hd__decap_3 PHY_11493 ();
 sky130_fd_sc_hd__decap_3 PHY_11494 ();
 sky130_fd_sc_hd__decap_3 PHY_11495 ();
 sky130_fd_sc_hd__decap_3 PHY_11496 ();
 sky130_fd_sc_hd__decap_3 PHY_11497 ();
 sky130_fd_sc_hd__decap_3 PHY_11498 ();
 sky130_fd_sc_hd__decap_3 PHY_11499 ();
 sky130_fd_sc_hd__decap_3 PHY_11500 ();
 sky130_fd_sc_hd__decap_3 PHY_11501 ();
 sky130_fd_sc_hd__decap_3 PHY_11502 ();
 sky130_fd_sc_hd__decap_3 PHY_11503 ();
 sky130_fd_sc_hd__decap_3 PHY_11504 ();
 sky130_fd_sc_hd__decap_3 PHY_11505 ();
 sky130_fd_sc_hd__decap_3 PHY_11506 ();
 sky130_fd_sc_hd__decap_3 PHY_11507 ();
 sky130_fd_sc_hd__decap_3 PHY_11508 ();
 sky130_fd_sc_hd__decap_3 PHY_11509 ();
 sky130_fd_sc_hd__decap_3 PHY_11510 ();
 sky130_fd_sc_hd__decap_3 PHY_11511 ();
 sky130_fd_sc_hd__decap_3 PHY_11512 ();
 sky130_fd_sc_hd__decap_3 PHY_11513 ();
 sky130_fd_sc_hd__decap_3 PHY_11514 ();
 sky130_fd_sc_hd__decap_3 PHY_11515 ();
 sky130_fd_sc_hd__decap_3 PHY_11516 ();
 sky130_fd_sc_hd__decap_3 PHY_11517 ();
 sky130_fd_sc_hd__decap_3 PHY_11518 ();
 sky130_fd_sc_hd__decap_3 PHY_11519 ();
 sky130_fd_sc_hd__decap_3 PHY_11520 ();
 sky130_fd_sc_hd__decap_3 PHY_11521 ();
 sky130_fd_sc_hd__decap_3 PHY_11522 ();
 sky130_fd_sc_hd__decap_3 PHY_11523 ();
 sky130_fd_sc_hd__decap_3 PHY_11524 ();
 sky130_fd_sc_hd__decap_3 PHY_11525 ();
 sky130_fd_sc_hd__decap_3 PHY_11526 ();
 sky130_fd_sc_hd__decap_3 PHY_11527 ();
 sky130_fd_sc_hd__decap_3 PHY_11528 ();
 sky130_fd_sc_hd__decap_3 PHY_11529 ();
 sky130_fd_sc_hd__decap_3 PHY_11530 ();
 sky130_fd_sc_hd__decap_3 PHY_11531 ();
 sky130_fd_sc_hd__decap_3 PHY_11532 ();
 sky130_fd_sc_hd__decap_3 PHY_11533 ();
 sky130_fd_sc_hd__decap_3 PHY_11534 ();
 sky130_fd_sc_hd__decap_3 PHY_11535 ();
 sky130_fd_sc_hd__decap_3 PHY_11536 ();
 sky130_fd_sc_hd__decap_3 PHY_11537 ();
 sky130_fd_sc_hd__decap_3 PHY_11538 ();
 sky130_fd_sc_hd__decap_3 PHY_11539 ();
 sky130_fd_sc_hd__decap_3 PHY_11540 ();
 sky130_fd_sc_hd__decap_3 PHY_11541 ();
 sky130_fd_sc_hd__decap_3 PHY_11542 ();
 sky130_fd_sc_hd__decap_3 PHY_11543 ();
 sky130_fd_sc_hd__decap_3 PHY_11544 ();
 sky130_fd_sc_hd__decap_3 PHY_11545 ();
 sky130_fd_sc_hd__decap_3 PHY_11546 ();
 sky130_fd_sc_hd__decap_3 PHY_11547 ();
 sky130_fd_sc_hd__decap_3 PHY_11548 ();
 sky130_fd_sc_hd__decap_3 PHY_11549 ();
 sky130_fd_sc_hd__decap_3 PHY_11550 ();
 sky130_fd_sc_hd__decap_3 PHY_11551 ();
 sky130_fd_sc_hd__decap_3 PHY_11552 ();
 sky130_fd_sc_hd__decap_3 PHY_11553 ();
 sky130_fd_sc_hd__decap_3 PHY_11554 ();
 sky130_fd_sc_hd__decap_3 PHY_11555 ();
 sky130_fd_sc_hd__decap_3 PHY_11556 ();
 sky130_fd_sc_hd__decap_3 PHY_11557 ();
 sky130_fd_sc_hd__decap_3 PHY_11558 ();
 sky130_fd_sc_hd__decap_3 PHY_11559 ();
 sky130_fd_sc_hd__decap_3 PHY_11560 ();
 sky130_fd_sc_hd__decap_3 PHY_11561 ();
 sky130_fd_sc_hd__decap_3 PHY_11562 ();
 sky130_fd_sc_hd__decap_3 PHY_11563 ();
 sky130_fd_sc_hd__decap_3 PHY_11564 ();
 sky130_fd_sc_hd__decap_3 PHY_11565 ();
 sky130_fd_sc_hd__decap_3 PHY_11566 ();
 sky130_fd_sc_hd__decap_3 PHY_11567 ();
 sky130_fd_sc_hd__decap_3 PHY_11568 ();
 sky130_fd_sc_hd__decap_3 PHY_11569 ();
 sky130_fd_sc_hd__decap_3 PHY_11570 ();
 sky130_fd_sc_hd__decap_3 PHY_11571 ();
 sky130_fd_sc_hd__decap_3 PHY_11572 ();
 sky130_fd_sc_hd__decap_3 PHY_11573 ();
 sky130_fd_sc_hd__decap_3 PHY_11574 ();
 sky130_fd_sc_hd__decap_3 PHY_11575 ();
 sky130_fd_sc_hd__decap_3 PHY_11576 ();
 sky130_fd_sc_hd__decap_3 PHY_11577 ();
 sky130_fd_sc_hd__decap_3 PHY_11578 ();
 sky130_fd_sc_hd__decap_3 PHY_11579 ();
 sky130_fd_sc_hd__decap_3 PHY_11580 ();
 sky130_fd_sc_hd__decap_3 PHY_11581 ();
 sky130_fd_sc_hd__decap_3 PHY_11582 ();
 sky130_fd_sc_hd__decap_3 PHY_11583 ();
 sky130_fd_sc_hd__decap_3 PHY_11584 ();
 sky130_fd_sc_hd__decap_3 PHY_11585 ();
 sky130_fd_sc_hd__decap_3 PHY_11586 ();
 sky130_fd_sc_hd__decap_3 PHY_11587 ();
 sky130_fd_sc_hd__decap_3 PHY_11588 ();
 sky130_fd_sc_hd__decap_3 PHY_11589 ();
 sky130_fd_sc_hd__decap_3 PHY_11590 ();
 sky130_fd_sc_hd__decap_3 PHY_11591 ();
 sky130_fd_sc_hd__decap_3 PHY_11592 ();
 sky130_fd_sc_hd__decap_3 PHY_11593 ();
 sky130_fd_sc_hd__decap_3 PHY_11594 ();
 sky130_fd_sc_hd__decap_3 PHY_11595 ();
 sky130_fd_sc_hd__decap_3 PHY_11596 ();
 sky130_fd_sc_hd__decap_3 PHY_11597 ();
 sky130_fd_sc_hd__decap_3 PHY_11598 ();
 sky130_fd_sc_hd__decap_3 PHY_11599 ();
 sky130_fd_sc_hd__decap_3 PHY_11600 ();
 sky130_fd_sc_hd__decap_3 PHY_11601 ();
 sky130_fd_sc_hd__decap_3 PHY_11602 ();
 sky130_fd_sc_hd__decap_3 PHY_11603 ();
 sky130_fd_sc_hd__decap_3 PHY_11604 ();
 sky130_fd_sc_hd__decap_3 PHY_11605 ();
 sky130_fd_sc_hd__decap_3 PHY_11606 ();
 sky130_fd_sc_hd__decap_3 PHY_11607 ();
 sky130_fd_sc_hd__decap_3 PHY_11608 ();
 sky130_fd_sc_hd__decap_3 PHY_11609 ();
 sky130_fd_sc_hd__decap_3 PHY_11610 ();
 sky130_fd_sc_hd__decap_3 PHY_11611 ();
 sky130_fd_sc_hd__decap_3 PHY_11612 ();
 sky130_fd_sc_hd__decap_3 PHY_11613 ();
 sky130_fd_sc_hd__decap_3 PHY_11614 ();
 sky130_fd_sc_hd__decap_3 PHY_11615 ();
 sky130_fd_sc_hd__decap_3 PHY_11616 ();
 sky130_fd_sc_hd__decap_3 PHY_11617 ();
 sky130_fd_sc_hd__decap_3 PHY_11618 ();
 sky130_fd_sc_hd__decap_3 PHY_11619 ();
 sky130_fd_sc_hd__decap_3 PHY_11620 ();
 sky130_fd_sc_hd__decap_3 PHY_11621 ();
 sky130_fd_sc_hd__decap_3 PHY_11622 ();
 sky130_fd_sc_hd__decap_3 PHY_11623 ();
 sky130_fd_sc_hd__decap_3 PHY_11624 ();
 sky130_fd_sc_hd__decap_3 PHY_11625 ();
 sky130_fd_sc_hd__decap_3 PHY_11626 ();
 sky130_fd_sc_hd__decap_3 PHY_11627 ();
 sky130_fd_sc_hd__decap_3 PHY_11628 ();
 sky130_fd_sc_hd__decap_3 PHY_11629 ();
 sky130_fd_sc_hd__decap_3 PHY_11630 ();
 sky130_fd_sc_hd__decap_3 PHY_11631 ();
 sky130_fd_sc_hd__decap_3 PHY_11632 ();
 sky130_fd_sc_hd__decap_3 PHY_11633 ();
 sky130_fd_sc_hd__decap_3 PHY_11634 ();
 sky130_fd_sc_hd__decap_3 PHY_11635 ();
 sky130_fd_sc_hd__decap_3 PHY_11636 ();
 sky130_fd_sc_hd__decap_3 PHY_11637 ();
 sky130_fd_sc_hd__decap_3 PHY_11638 ();
 sky130_fd_sc_hd__decap_3 PHY_11639 ();
 sky130_fd_sc_hd__decap_3 PHY_11640 ();
 sky130_fd_sc_hd__decap_3 PHY_11641 ();
 sky130_fd_sc_hd__decap_3 PHY_11642 ();
 sky130_fd_sc_hd__decap_3 PHY_11643 ();
 sky130_fd_sc_hd__decap_3 PHY_11644 ();
 sky130_fd_sc_hd__decap_3 PHY_11645 ();
 sky130_fd_sc_hd__decap_3 PHY_11646 ();
 sky130_fd_sc_hd__decap_3 PHY_11647 ();
 sky130_fd_sc_hd__decap_3 PHY_11648 ();
 sky130_fd_sc_hd__decap_3 PHY_11649 ();
 sky130_fd_sc_hd__decap_3 PHY_11650 ();
 sky130_fd_sc_hd__decap_3 PHY_11651 ();
 sky130_fd_sc_hd__decap_3 PHY_11652 ();
 sky130_fd_sc_hd__decap_3 PHY_11653 ();
 sky130_fd_sc_hd__decap_3 PHY_11654 ();
 sky130_fd_sc_hd__decap_3 PHY_11655 ();
 sky130_fd_sc_hd__decap_3 PHY_11656 ();
 sky130_fd_sc_hd__decap_3 PHY_11657 ();
 sky130_fd_sc_hd__decap_3 PHY_11658 ();
 sky130_fd_sc_hd__decap_3 PHY_11659 ();
 sky130_fd_sc_hd__decap_3 PHY_11660 ();
 sky130_fd_sc_hd__decap_3 PHY_11661 ();
 sky130_fd_sc_hd__decap_3 PHY_11662 ();
 sky130_fd_sc_hd__decap_3 PHY_11663 ();
 sky130_fd_sc_hd__decap_3 PHY_11664 ();
 sky130_fd_sc_hd__decap_3 PHY_11665 ();
 sky130_fd_sc_hd__decap_3 PHY_11666 ();
 sky130_fd_sc_hd__decap_3 PHY_11667 ();
 sky130_fd_sc_hd__decap_3 PHY_11668 ();
 sky130_fd_sc_hd__decap_3 PHY_11669 ();
 sky130_fd_sc_hd__decap_3 PHY_11670 ();
 sky130_fd_sc_hd__decap_3 PHY_11671 ();
 sky130_fd_sc_hd__decap_3 PHY_11672 ();
 sky130_fd_sc_hd__decap_3 PHY_11673 ();
 sky130_fd_sc_hd__decap_3 PHY_11674 ();
 sky130_fd_sc_hd__decap_3 PHY_11675 ();
 sky130_fd_sc_hd__decap_3 PHY_11676 ();
 sky130_fd_sc_hd__decap_3 PHY_11677 ();
 sky130_fd_sc_hd__decap_3 PHY_11678 ();
 sky130_fd_sc_hd__decap_3 PHY_11679 ();
 sky130_fd_sc_hd__decap_3 PHY_11680 ();
 sky130_fd_sc_hd__decap_3 PHY_11681 ();
 sky130_fd_sc_hd__decap_3 PHY_11682 ();
 sky130_fd_sc_hd__decap_3 PHY_11683 ();
 sky130_fd_sc_hd__decap_3 PHY_11684 ();
 sky130_fd_sc_hd__decap_3 PHY_11685 ();
 sky130_fd_sc_hd__decap_3 PHY_11686 ();
 sky130_fd_sc_hd__decap_3 PHY_11687 ();
 sky130_fd_sc_hd__decap_3 PHY_11688 ();
 sky130_fd_sc_hd__decap_3 PHY_11689 ();
 sky130_fd_sc_hd__decap_3 PHY_11690 ();
 sky130_fd_sc_hd__decap_3 PHY_11691 ();
 sky130_fd_sc_hd__decap_3 PHY_11692 ();
 sky130_fd_sc_hd__decap_3 PHY_11693 ();
 sky130_fd_sc_hd__decap_3 PHY_11694 ();
 sky130_fd_sc_hd__decap_3 PHY_11695 ();
 sky130_fd_sc_hd__decap_3 PHY_11696 ();
 sky130_fd_sc_hd__decap_3 PHY_11697 ();
 sky130_fd_sc_hd__decap_3 PHY_11698 ();
 sky130_fd_sc_hd__decap_3 PHY_11699 ();
 sky130_fd_sc_hd__decap_3 PHY_11700 ();
 sky130_fd_sc_hd__decap_3 PHY_11701 ();
 sky130_fd_sc_hd__decap_3 PHY_11702 ();
 sky130_fd_sc_hd__decap_3 PHY_11703 ();
 sky130_fd_sc_hd__decap_3 PHY_11704 ();
 sky130_fd_sc_hd__decap_3 PHY_11705 ();
 sky130_fd_sc_hd__decap_3 PHY_11706 ();
 sky130_fd_sc_hd__decap_3 PHY_11707 ();
 sky130_fd_sc_hd__decap_3 PHY_11708 ();
 sky130_fd_sc_hd__decap_3 PHY_11709 ();
 sky130_fd_sc_hd__decap_3 PHY_11710 ();
 sky130_fd_sc_hd__decap_3 PHY_11711 ();
 sky130_fd_sc_hd__decap_3 PHY_11712 ();
 sky130_fd_sc_hd__decap_3 PHY_11713 ();
 sky130_fd_sc_hd__decap_3 PHY_11714 ();
 sky130_fd_sc_hd__decap_3 PHY_11715 ();
 sky130_fd_sc_hd__decap_3 PHY_11716 ();
 sky130_fd_sc_hd__decap_3 PHY_11717 ();
 sky130_fd_sc_hd__decap_3 PHY_11718 ();
 sky130_fd_sc_hd__decap_3 PHY_11719 ();
 sky130_fd_sc_hd__decap_3 PHY_11720 ();
 sky130_fd_sc_hd__decap_3 PHY_11721 ();
 sky130_fd_sc_hd__decap_3 PHY_11722 ();
 sky130_fd_sc_hd__decap_3 PHY_11723 ();
 sky130_fd_sc_hd__decap_3 PHY_11724 ();
 sky130_fd_sc_hd__decap_3 PHY_11725 ();
 sky130_fd_sc_hd__decap_3 PHY_11726 ();
 sky130_fd_sc_hd__decap_3 PHY_11727 ();
 sky130_fd_sc_hd__decap_3 PHY_11728 ();
 sky130_fd_sc_hd__decap_3 PHY_11729 ();
 sky130_fd_sc_hd__decap_3 PHY_11730 ();
 sky130_fd_sc_hd__decap_3 PHY_11731 ();
 sky130_fd_sc_hd__decap_3 PHY_11732 ();
 sky130_fd_sc_hd__decap_3 PHY_11733 ();
 sky130_fd_sc_hd__decap_3 PHY_11734 ();
 sky130_fd_sc_hd__decap_3 PHY_11735 ();
 sky130_fd_sc_hd__decap_3 PHY_11736 ();
 sky130_fd_sc_hd__decap_3 PHY_11737 ();
 sky130_fd_sc_hd__decap_3 PHY_11738 ();
 sky130_fd_sc_hd__decap_3 PHY_11739 ();
 sky130_fd_sc_hd__decap_3 PHY_11740 ();
 sky130_fd_sc_hd__decap_3 PHY_11741 ();
 sky130_fd_sc_hd__decap_3 PHY_11742 ();
 sky130_fd_sc_hd__decap_3 PHY_11743 ();
 sky130_fd_sc_hd__decap_3 PHY_11744 ();
 sky130_fd_sc_hd__decap_3 PHY_11745 ();
 sky130_fd_sc_hd__decap_3 PHY_11746 ();
 sky130_fd_sc_hd__decap_3 PHY_11747 ();
 sky130_fd_sc_hd__decap_3 PHY_11748 ();
 sky130_fd_sc_hd__decap_3 PHY_11749 ();
 sky130_fd_sc_hd__decap_3 PHY_11750 ();
 sky130_fd_sc_hd__decap_3 PHY_11751 ();
 sky130_fd_sc_hd__decap_3 PHY_11752 ();
 sky130_fd_sc_hd__decap_3 PHY_11753 ();
 sky130_fd_sc_hd__decap_3 PHY_11754 ();
 sky130_fd_sc_hd__decap_3 PHY_11755 ();
 sky130_fd_sc_hd__decap_3 PHY_11756 ();
 sky130_fd_sc_hd__decap_3 PHY_11757 ();
 sky130_fd_sc_hd__decap_3 PHY_11758 ();
 sky130_fd_sc_hd__decap_3 PHY_11759 ();
 sky130_fd_sc_hd__decap_3 PHY_11760 ();
 sky130_fd_sc_hd__decap_3 PHY_11761 ();
 sky130_fd_sc_hd__decap_3 PHY_11762 ();
 sky130_fd_sc_hd__decap_3 PHY_11763 ();
 sky130_fd_sc_hd__decap_3 PHY_11764 ();
 sky130_fd_sc_hd__decap_3 PHY_11765 ();
 sky130_fd_sc_hd__decap_3 PHY_11766 ();
 sky130_fd_sc_hd__decap_3 PHY_11767 ();
 sky130_fd_sc_hd__decap_3 PHY_11768 ();
 sky130_fd_sc_hd__decap_3 PHY_11769 ();
 sky130_fd_sc_hd__decap_3 PHY_11770 ();
 sky130_fd_sc_hd__decap_3 PHY_11771 ();
 sky130_fd_sc_hd__decap_3 PHY_11772 ();
 sky130_fd_sc_hd__decap_3 PHY_11773 ();
 sky130_fd_sc_hd__decap_3 PHY_11774 ();
 sky130_fd_sc_hd__decap_3 PHY_11775 ();
 sky130_fd_sc_hd__decap_3 PHY_11776 ();
 sky130_fd_sc_hd__decap_3 PHY_11777 ();
 sky130_fd_sc_hd__decap_3 PHY_11778 ();
 sky130_fd_sc_hd__decap_3 PHY_11779 ();
 sky130_fd_sc_hd__decap_3 PHY_11780 ();
 sky130_fd_sc_hd__decap_3 PHY_11781 ();
 sky130_fd_sc_hd__decap_3 PHY_11782 ();
 sky130_fd_sc_hd__decap_3 PHY_11783 ();
 sky130_fd_sc_hd__decap_3 PHY_11784 ();
 sky130_fd_sc_hd__decap_3 PHY_11785 ();
 sky130_fd_sc_hd__decap_3 PHY_11786 ();
 sky130_fd_sc_hd__decap_3 PHY_11787 ();
 sky130_fd_sc_hd__decap_3 PHY_11788 ();
 sky130_fd_sc_hd__decap_3 PHY_11789 ();
 sky130_fd_sc_hd__decap_3 PHY_11790 ();
 sky130_fd_sc_hd__decap_3 PHY_11791 ();
 sky130_fd_sc_hd__decap_3 PHY_11792 ();
 sky130_fd_sc_hd__decap_3 PHY_11793 ();
 sky130_fd_sc_hd__decap_3 PHY_11794 ();
 sky130_fd_sc_hd__decap_3 PHY_11795 ();
 sky130_fd_sc_hd__decap_3 PHY_11796 ();
 sky130_fd_sc_hd__decap_3 PHY_11797 ();
 sky130_fd_sc_hd__decap_3 PHY_11798 ();
 sky130_fd_sc_hd__decap_3 PHY_11799 ();
 sky130_fd_sc_hd__decap_3 PHY_11800 ();
 sky130_fd_sc_hd__decap_3 PHY_11801 ();
 sky130_fd_sc_hd__decap_3 PHY_11802 ();
 sky130_fd_sc_hd__decap_3 PHY_11803 ();
 sky130_fd_sc_hd__decap_3 PHY_11804 ();
 sky130_fd_sc_hd__decap_3 PHY_11805 ();
 sky130_fd_sc_hd__decap_3 PHY_11806 ();
 sky130_fd_sc_hd__decap_3 PHY_11807 ();
 sky130_fd_sc_hd__decap_3 PHY_11808 ();
 sky130_fd_sc_hd__decap_3 PHY_11809 ();
 sky130_fd_sc_hd__decap_3 PHY_11810 ();
 sky130_fd_sc_hd__decap_3 PHY_11811 ();
 sky130_fd_sc_hd__decap_3 PHY_11812 ();
 sky130_fd_sc_hd__decap_3 PHY_11813 ();
 sky130_fd_sc_hd__decap_3 PHY_11814 ();
 sky130_fd_sc_hd__decap_3 PHY_11815 ();
 sky130_fd_sc_hd__decap_3 PHY_11816 ();
 sky130_fd_sc_hd__decap_3 PHY_11817 ();
 sky130_fd_sc_hd__decap_3 PHY_11818 ();
 sky130_fd_sc_hd__decap_3 PHY_11819 ();
 sky130_fd_sc_hd__decap_3 PHY_11820 ();
 sky130_fd_sc_hd__decap_3 PHY_11821 ();
 sky130_fd_sc_hd__decap_3 PHY_11822 ();
 sky130_fd_sc_hd__decap_3 PHY_11823 ();
 sky130_fd_sc_hd__decap_3 PHY_11824 ();
 sky130_fd_sc_hd__decap_3 PHY_11825 ();
 sky130_fd_sc_hd__decap_3 PHY_11826 ();
 sky130_fd_sc_hd__decap_3 PHY_11827 ();
 sky130_fd_sc_hd__decap_3 PHY_11828 ();
 sky130_fd_sc_hd__decap_3 PHY_11829 ();
 sky130_fd_sc_hd__decap_3 PHY_11830 ();
 sky130_fd_sc_hd__decap_3 PHY_11831 ();
 sky130_fd_sc_hd__decap_3 PHY_11832 ();
 sky130_fd_sc_hd__decap_3 PHY_11833 ();
 sky130_fd_sc_hd__decap_3 PHY_11834 ();
 sky130_fd_sc_hd__decap_3 PHY_11835 ();
 sky130_fd_sc_hd__decap_3 PHY_11836 ();
 sky130_fd_sc_hd__decap_3 PHY_11837 ();
 sky130_fd_sc_hd__decap_3 PHY_11838 ();
 sky130_fd_sc_hd__decap_3 PHY_11839 ();
 sky130_fd_sc_hd__decap_3 PHY_11840 ();
 sky130_fd_sc_hd__decap_3 PHY_11841 ();
 sky130_fd_sc_hd__decap_3 PHY_11842 ();
 sky130_fd_sc_hd__decap_3 PHY_11843 ();
 sky130_fd_sc_hd__decap_3 PHY_11844 ();
 sky130_fd_sc_hd__decap_3 PHY_11845 ();
 sky130_fd_sc_hd__decap_3 PHY_11846 ();
 sky130_fd_sc_hd__decap_3 PHY_11847 ();
 sky130_fd_sc_hd__decap_3 PHY_11848 ();
 sky130_fd_sc_hd__decap_3 PHY_11849 ();
 sky130_fd_sc_hd__decap_3 PHY_11850 ();
 sky130_fd_sc_hd__decap_3 PHY_11851 ();
 sky130_fd_sc_hd__decap_3 PHY_11852 ();
 sky130_fd_sc_hd__decap_3 PHY_11853 ();
 sky130_fd_sc_hd__decap_3 PHY_11854 ();
 sky130_fd_sc_hd__decap_3 PHY_11855 ();
 sky130_fd_sc_hd__decap_3 PHY_11856 ();
 sky130_fd_sc_hd__decap_3 PHY_11857 ();
 sky130_fd_sc_hd__decap_3 PHY_11858 ();
 sky130_fd_sc_hd__decap_3 PHY_11859 ();
 sky130_fd_sc_hd__decap_3 PHY_11860 ();
 sky130_fd_sc_hd__decap_3 PHY_11861 ();
 sky130_fd_sc_hd__decap_3 PHY_11862 ();
 sky130_fd_sc_hd__decap_3 PHY_11863 ();
 sky130_fd_sc_hd__decap_3 PHY_11864 ();
 sky130_fd_sc_hd__decap_3 PHY_11865 ();
 sky130_fd_sc_hd__decap_3 PHY_11866 ();
 sky130_fd_sc_hd__decap_3 PHY_11867 ();
 sky130_fd_sc_hd__decap_3 PHY_11868 ();
 sky130_fd_sc_hd__decap_3 PHY_11869 ();
 sky130_fd_sc_hd__decap_3 PHY_11870 ();
 sky130_fd_sc_hd__decap_3 PHY_11871 ();
 sky130_fd_sc_hd__decap_3 PHY_11872 ();
 sky130_fd_sc_hd__decap_3 PHY_11873 ();
 sky130_fd_sc_hd__decap_3 PHY_11874 ();
 sky130_fd_sc_hd__decap_3 PHY_11875 ();
 sky130_fd_sc_hd__decap_3 PHY_11876 ();
 sky130_fd_sc_hd__decap_3 PHY_11877 ();
 sky130_fd_sc_hd__decap_3 PHY_11878 ();
 sky130_fd_sc_hd__decap_3 PHY_11879 ();
 sky130_fd_sc_hd__decap_3 PHY_11880 ();
 sky130_fd_sc_hd__decap_3 PHY_11881 ();
 sky130_fd_sc_hd__decap_3 PHY_11882 ();
 sky130_fd_sc_hd__decap_3 PHY_11883 ();
 sky130_fd_sc_hd__decap_3 PHY_11884 ();
 sky130_fd_sc_hd__decap_3 PHY_11885 ();
 sky130_fd_sc_hd__decap_3 PHY_11886 ();
 sky130_fd_sc_hd__decap_3 PHY_11887 ();
 sky130_fd_sc_hd__decap_3 PHY_11888 ();
 sky130_fd_sc_hd__decap_3 PHY_11889 ();
 sky130_fd_sc_hd__decap_3 PHY_11890 ();
 sky130_fd_sc_hd__decap_3 PHY_11891 ();
 sky130_fd_sc_hd__decap_3 PHY_11892 ();
 sky130_fd_sc_hd__decap_3 PHY_11893 ();
 sky130_fd_sc_hd__decap_3 PHY_11894 ();
 sky130_fd_sc_hd__decap_3 PHY_11895 ();
 sky130_fd_sc_hd__decap_3 PHY_11896 ();
 sky130_fd_sc_hd__decap_3 PHY_11897 ();
 sky130_fd_sc_hd__decap_3 PHY_11898 ();
 sky130_fd_sc_hd__decap_3 PHY_11899 ();
 sky130_fd_sc_hd__decap_3 PHY_11900 ();
 sky130_fd_sc_hd__decap_3 PHY_11901 ();
 sky130_fd_sc_hd__decap_3 PHY_11902 ();
 sky130_fd_sc_hd__decap_3 PHY_11903 ();
 sky130_fd_sc_hd__decap_3 PHY_11904 ();
 sky130_fd_sc_hd__decap_3 PHY_11905 ();
 sky130_fd_sc_hd__decap_3 PHY_11906 ();
 sky130_fd_sc_hd__decap_3 PHY_11907 ();
 sky130_fd_sc_hd__decap_3 PHY_11908 ();
 sky130_fd_sc_hd__decap_3 PHY_11909 ();
 sky130_fd_sc_hd__decap_3 PHY_11910 ();
 sky130_fd_sc_hd__decap_3 PHY_11911 ();
 sky130_fd_sc_hd__decap_3 PHY_11912 ();
 sky130_fd_sc_hd__decap_3 PHY_11913 ();
 sky130_fd_sc_hd__decap_3 PHY_11914 ();
 sky130_fd_sc_hd__decap_3 PHY_11915 ();
 sky130_fd_sc_hd__decap_3 PHY_11916 ();
 sky130_fd_sc_hd__decap_3 PHY_11917 ();
 sky130_fd_sc_hd__decap_3 PHY_11918 ();
 sky130_fd_sc_hd__decap_3 PHY_11919 ();
 sky130_fd_sc_hd__decap_3 PHY_11920 ();
 sky130_fd_sc_hd__decap_3 PHY_11921 ();
 sky130_fd_sc_hd__decap_3 PHY_11922 ();
 sky130_fd_sc_hd__decap_3 PHY_11923 ();
 sky130_fd_sc_hd__decap_3 PHY_11924 ();
 sky130_fd_sc_hd__decap_3 PHY_11925 ();
 sky130_fd_sc_hd__decap_3 PHY_11926 ();
 sky130_fd_sc_hd__decap_3 PHY_11927 ();
 sky130_fd_sc_hd__decap_3 PHY_11928 ();
 sky130_fd_sc_hd__decap_3 PHY_11929 ();
 sky130_fd_sc_hd__decap_3 PHY_11930 ();
 sky130_fd_sc_hd__decap_3 PHY_11931 ();
 sky130_fd_sc_hd__decap_3 PHY_11932 ();
 sky130_fd_sc_hd__decap_3 PHY_11933 ();
 sky130_fd_sc_hd__decap_3 PHY_11934 ();
 sky130_fd_sc_hd__decap_3 PHY_11935 ();
 sky130_fd_sc_hd__decap_3 PHY_11936 ();
 sky130_fd_sc_hd__decap_3 PHY_11937 ();
 sky130_fd_sc_hd__decap_3 PHY_11938 ();
 sky130_fd_sc_hd__decap_3 PHY_11939 ();
 sky130_fd_sc_hd__decap_3 PHY_11940 ();
 sky130_fd_sc_hd__decap_3 PHY_11941 ();
 sky130_fd_sc_hd__decap_3 PHY_11942 ();
 sky130_fd_sc_hd__decap_3 PHY_11943 ();
 sky130_fd_sc_hd__decap_3 PHY_11944 ();
 sky130_fd_sc_hd__decap_3 PHY_11945 ();
 sky130_fd_sc_hd__decap_3 PHY_11946 ();
 sky130_fd_sc_hd__decap_3 PHY_11947 ();
 sky130_fd_sc_hd__decap_3 PHY_11948 ();
 sky130_fd_sc_hd__decap_3 PHY_11949 ();
 sky130_fd_sc_hd__decap_3 PHY_11950 ();
 sky130_fd_sc_hd__decap_3 PHY_11951 ();
 sky130_fd_sc_hd__decap_3 PHY_11952 ();
 sky130_fd_sc_hd__decap_3 PHY_11953 ();
 sky130_fd_sc_hd__decap_3 PHY_11954 ();
 sky130_fd_sc_hd__decap_3 PHY_11955 ();
 sky130_fd_sc_hd__decap_3 PHY_11956 ();
 sky130_fd_sc_hd__decap_3 PHY_11957 ();
 sky130_fd_sc_hd__decap_3 PHY_11958 ();
 sky130_fd_sc_hd__decap_3 PHY_11959 ();
 sky130_fd_sc_hd__decap_3 PHY_11960 ();
 sky130_fd_sc_hd__decap_3 PHY_11961 ();
 sky130_fd_sc_hd__decap_3 PHY_11962 ();
 sky130_fd_sc_hd__decap_3 PHY_11963 ();
 sky130_fd_sc_hd__decap_3 PHY_11964 ();
 sky130_fd_sc_hd__decap_3 PHY_11965 ();
 sky130_fd_sc_hd__decap_3 PHY_11966 ();
 sky130_fd_sc_hd__decap_3 PHY_11967 ();
 sky130_fd_sc_hd__decap_3 PHY_11968 ();
 sky130_fd_sc_hd__decap_3 PHY_11969 ();
 sky130_fd_sc_hd__decap_3 PHY_11970 ();
 sky130_fd_sc_hd__decap_3 PHY_11971 ();
 sky130_fd_sc_hd__decap_3 PHY_11972 ();
 sky130_fd_sc_hd__decap_3 PHY_11973 ();
 sky130_fd_sc_hd__decap_3 PHY_11974 ();
 sky130_fd_sc_hd__decap_3 PHY_11975 ();
 sky130_fd_sc_hd__decap_3 PHY_11976 ();
 sky130_fd_sc_hd__decap_3 PHY_11977 ();
 sky130_fd_sc_hd__decap_3 PHY_11978 ();
 sky130_fd_sc_hd__decap_3 PHY_11979 ();
 sky130_fd_sc_hd__decap_3 PHY_11980 ();
 sky130_fd_sc_hd__decap_3 PHY_11981 ();
 sky130_fd_sc_hd__decap_3 PHY_11982 ();
 sky130_fd_sc_hd__decap_3 PHY_11983 ();
 sky130_fd_sc_hd__decap_3 PHY_11984 ();
 sky130_fd_sc_hd__decap_3 PHY_11985 ();
 sky130_fd_sc_hd__decap_3 PHY_11986 ();
 sky130_fd_sc_hd__decap_3 PHY_11987 ();
 sky130_fd_sc_hd__decap_3 PHY_11988 ();
 sky130_fd_sc_hd__decap_3 PHY_11989 ();
 sky130_fd_sc_hd__decap_3 PHY_11990 ();
 sky130_fd_sc_hd__decap_3 PHY_11991 ();
 sky130_fd_sc_hd__decap_3 PHY_11992 ();
 sky130_fd_sc_hd__decap_3 PHY_11993 ();
 sky130_fd_sc_hd__decap_3 PHY_11994 ();
 sky130_fd_sc_hd__decap_3 PHY_11995 ();
 sky130_fd_sc_hd__decap_3 PHY_11996 ();
 sky130_fd_sc_hd__decap_3 PHY_11997 ();
 sky130_fd_sc_hd__decap_3 PHY_11998 ();
 sky130_fd_sc_hd__decap_3 PHY_11999 ();
 sky130_fd_sc_hd__decap_3 PHY_12000 ();
 sky130_fd_sc_hd__decap_3 PHY_12001 ();
 sky130_fd_sc_hd__decap_3 PHY_12002 ();
 sky130_fd_sc_hd__decap_3 PHY_12003 ();
 sky130_fd_sc_hd__decap_3 PHY_12004 ();
 sky130_fd_sc_hd__decap_3 PHY_12005 ();
 sky130_fd_sc_hd__decap_3 PHY_12006 ();
 sky130_fd_sc_hd__decap_3 PHY_12007 ();
 sky130_fd_sc_hd__decap_3 PHY_12008 ();
 sky130_fd_sc_hd__decap_3 PHY_12009 ();
 sky130_fd_sc_hd__decap_3 PHY_12010 ();
 sky130_fd_sc_hd__decap_3 PHY_12011 ();
 sky130_fd_sc_hd__decap_3 PHY_12012 ();
 sky130_fd_sc_hd__decap_3 PHY_12013 ();
 sky130_fd_sc_hd__decap_3 PHY_12014 ();
 sky130_fd_sc_hd__decap_3 PHY_12015 ();
 sky130_fd_sc_hd__decap_3 PHY_12016 ();
 sky130_fd_sc_hd__decap_3 PHY_12017 ();
 sky130_fd_sc_hd__decap_3 PHY_12018 ();
 sky130_fd_sc_hd__decap_3 PHY_12019 ();
 sky130_fd_sc_hd__decap_3 PHY_12020 ();
 sky130_fd_sc_hd__decap_3 PHY_12021 ();
 sky130_fd_sc_hd__decap_3 PHY_12022 ();
 sky130_fd_sc_hd__decap_3 PHY_12023 ();
 sky130_fd_sc_hd__decap_3 PHY_12024 ();
 sky130_fd_sc_hd__decap_3 PHY_12025 ();
 sky130_fd_sc_hd__decap_3 PHY_12026 ();
 sky130_fd_sc_hd__decap_3 PHY_12027 ();
 sky130_fd_sc_hd__decap_3 PHY_12028 ();
 sky130_fd_sc_hd__decap_3 PHY_12029 ();
 sky130_fd_sc_hd__decap_3 PHY_12030 ();
 sky130_fd_sc_hd__decap_3 PHY_12031 ();
 sky130_fd_sc_hd__decap_3 PHY_12032 ();
 sky130_fd_sc_hd__decap_3 PHY_12033 ();
 sky130_fd_sc_hd__decap_3 PHY_12034 ();
 sky130_fd_sc_hd__decap_3 PHY_12035 ();
 sky130_fd_sc_hd__decap_3 PHY_12036 ();
 sky130_fd_sc_hd__decap_3 PHY_12037 ();
 sky130_fd_sc_hd__decap_3 PHY_12038 ();
 sky130_fd_sc_hd__decap_3 PHY_12039 ();
 sky130_fd_sc_hd__decap_3 PHY_12040 ();
 sky130_fd_sc_hd__decap_3 PHY_12041 ();
 sky130_fd_sc_hd__decap_3 PHY_12042 ();
 sky130_fd_sc_hd__decap_3 PHY_12043 ();
 sky130_fd_sc_hd__decap_3 PHY_12044 ();
 sky130_fd_sc_hd__decap_3 PHY_12045 ();
 sky130_fd_sc_hd__decap_3 PHY_12046 ();
 sky130_fd_sc_hd__decap_3 PHY_12047 ();
 sky130_fd_sc_hd__decap_3 PHY_12048 ();
 sky130_fd_sc_hd__decap_3 PHY_12049 ();
 sky130_fd_sc_hd__decap_3 PHY_12050 ();
 sky130_fd_sc_hd__decap_3 PHY_12051 ();
 sky130_fd_sc_hd__decap_3 PHY_12052 ();
 sky130_fd_sc_hd__decap_3 PHY_12053 ();
 sky130_fd_sc_hd__decap_3 PHY_12054 ();
 sky130_fd_sc_hd__decap_3 PHY_12055 ();
 sky130_fd_sc_hd__decap_3 PHY_12056 ();
 sky130_fd_sc_hd__decap_3 PHY_12057 ();
 sky130_fd_sc_hd__decap_3 PHY_12058 ();
 sky130_fd_sc_hd__decap_3 PHY_12059 ();
 sky130_fd_sc_hd__decap_3 PHY_12060 ();
 sky130_fd_sc_hd__decap_3 PHY_12061 ();
 sky130_fd_sc_hd__decap_3 PHY_12062 ();
 sky130_fd_sc_hd__decap_3 PHY_12063 ();
 sky130_fd_sc_hd__decap_3 PHY_12064 ();
 sky130_fd_sc_hd__decap_3 PHY_12065 ();
 sky130_fd_sc_hd__decap_3 PHY_12066 ();
 sky130_fd_sc_hd__decap_3 PHY_12067 ();
 sky130_fd_sc_hd__decap_3 PHY_12068 ();
 sky130_fd_sc_hd__decap_3 PHY_12069 ();
 sky130_fd_sc_hd__decap_3 PHY_12070 ();
 sky130_fd_sc_hd__decap_3 PHY_12071 ();
 sky130_fd_sc_hd__decap_3 PHY_12072 ();
 sky130_fd_sc_hd__decap_3 PHY_12073 ();
 sky130_fd_sc_hd__decap_3 PHY_12074 ();
 sky130_fd_sc_hd__decap_3 PHY_12075 ();
 sky130_fd_sc_hd__decap_3 PHY_12076 ();
 sky130_fd_sc_hd__decap_3 PHY_12077 ();
 sky130_fd_sc_hd__decap_3 PHY_12078 ();
 sky130_fd_sc_hd__decap_3 PHY_12079 ();
 sky130_fd_sc_hd__decap_3 PHY_12080 ();
 sky130_fd_sc_hd__decap_3 PHY_12081 ();
 sky130_fd_sc_hd__decap_3 PHY_12082 ();
 sky130_fd_sc_hd__decap_3 PHY_12083 ();
 sky130_fd_sc_hd__decap_3 PHY_12084 ();
 sky130_fd_sc_hd__decap_3 PHY_12085 ();
 sky130_fd_sc_hd__decap_3 PHY_12086 ();
 sky130_fd_sc_hd__decap_3 PHY_12087 ();
 sky130_fd_sc_hd__decap_3 PHY_12088 ();
 sky130_fd_sc_hd__decap_3 PHY_12089 ();
 sky130_fd_sc_hd__decap_3 PHY_12090 ();
 sky130_fd_sc_hd__decap_3 PHY_12091 ();
 sky130_fd_sc_hd__decap_3 PHY_12092 ();
 sky130_fd_sc_hd__decap_3 PHY_12093 ();
 sky130_fd_sc_hd__decap_3 PHY_12094 ();
 sky130_fd_sc_hd__decap_3 PHY_12095 ();
 sky130_fd_sc_hd__decap_3 PHY_12096 ();
 sky130_fd_sc_hd__decap_3 PHY_12097 ();
 sky130_fd_sc_hd__decap_3 PHY_12098 ();
 sky130_fd_sc_hd__decap_3 PHY_12099 ();
 sky130_fd_sc_hd__decap_3 PHY_12100 ();
 sky130_fd_sc_hd__decap_3 PHY_12101 ();
 sky130_fd_sc_hd__decap_3 PHY_12102 ();
 sky130_fd_sc_hd__decap_3 PHY_12103 ();
 sky130_fd_sc_hd__decap_3 PHY_12104 ();
 sky130_fd_sc_hd__decap_3 PHY_12105 ();
 sky130_fd_sc_hd__decap_3 PHY_12106 ();
 sky130_fd_sc_hd__decap_3 PHY_12107 ();
 sky130_fd_sc_hd__decap_3 PHY_12108 ();
 sky130_fd_sc_hd__decap_3 PHY_12109 ();
 sky130_fd_sc_hd__decap_3 PHY_12110 ();
 sky130_fd_sc_hd__decap_3 PHY_12111 ();
 sky130_fd_sc_hd__decap_3 PHY_12112 ();
 sky130_fd_sc_hd__decap_3 PHY_12113 ();
 sky130_fd_sc_hd__decap_3 PHY_12114 ();
 sky130_fd_sc_hd__decap_3 PHY_12115 ();
 sky130_fd_sc_hd__decap_3 PHY_12116 ();
 sky130_fd_sc_hd__decap_3 PHY_12117 ();
 sky130_fd_sc_hd__decap_3 PHY_12118 ();
 sky130_fd_sc_hd__decap_3 PHY_12119 ();
 sky130_fd_sc_hd__decap_3 PHY_12120 ();
 sky130_fd_sc_hd__decap_3 PHY_12121 ();
 sky130_fd_sc_hd__decap_3 PHY_12122 ();
 sky130_fd_sc_hd__decap_3 PHY_12123 ();
 sky130_fd_sc_hd__decap_3 PHY_12124 ();
 sky130_fd_sc_hd__decap_3 PHY_12125 ();
 sky130_fd_sc_hd__decap_3 PHY_12126 ();
 sky130_fd_sc_hd__decap_3 PHY_12127 ();
 sky130_fd_sc_hd__decap_3 PHY_12128 ();
 sky130_fd_sc_hd__decap_3 PHY_12129 ();
 sky130_fd_sc_hd__decap_3 PHY_12130 ();
 sky130_fd_sc_hd__decap_3 PHY_12131 ();
 sky130_fd_sc_hd__decap_3 PHY_12132 ();
 sky130_fd_sc_hd__decap_3 PHY_12133 ();
 sky130_fd_sc_hd__decap_3 PHY_12134 ();
 sky130_fd_sc_hd__decap_3 PHY_12135 ();
 sky130_fd_sc_hd__decap_3 PHY_12136 ();
 sky130_fd_sc_hd__decap_3 PHY_12137 ();
 sky130_fd_sc_hd__decap_3 PHY_12138 ();
 sky130_fd_sc_hd__decap_3 PHY_12139 ();
 sky130_fd_sc_hd__decap_3 PHY_12140 ();
 sky130_fd_sc_hd__decap_3 PHY_12141 ();
 sky130_fd_sc_hd__decap_3 PHY_12142 ();
 sky130_fd_sc_hd__decap_3 PHY_12143 ();
 sky130_fd_sc_hd__decap_3 PHY_12144 ();
 sky130_fd_sc_hd__decap_3 PHY_12145 ();
 sky130_fd_sc_hd__decap_3 PHY_12146 ();
 sky130_fd_sc_hd__decap_3 PHY_12147 ();
 sky130_fd_sc_hd__decap_3 PHY_12148 ();
 sky130_fd_sc_hd__decap_3 PHY_12149 ();
 sky130_fd_sc_hd__decap_3 PHY_12150 ();
 sky130_fd_sc_hd__decap_3 PHY_12151 ();
 sky130_fd_sc_hd__decap_3 PHY_12152 ();
 sky130_fd_sc_hd__decap_3 PHY_12153 ();
 sky130_fd_sc_hd__decap_3 PHY_12154 ();
 sky130_fd_sc_hd__decap_3 PHY_12155 ();
 sky130_fd_sc_hd__decap_3 PHY_12156 ();
 sky130_fd_sc_hd__decap_3 PHY_12157 ();
 sky130_fd_sc_hd__decap_3 PHY_12158 ();
 sky130_fd_sc_hd__decap_3 PHY_12159 ();
 sky130_fd_sc_hd__decap_3 PHY_12160 ();
 sky130_fd_sc_hd__decap_3 PHY_12161 ();
 sky130_fd_sc_hd__decap_3 PHY_12162 ();
 sky130_fd_sc_hd__decap_3 PHY_12163 ();
 sky130_fd_sc_hd__decap_3 PHY_12164 ();
 sky130_fd_sc_hd__decap_3 PHY_12165 ();
 sky130_fd_sc_hd__decap_3 PHY_12166 ();
 sky130_fd_sc_hd__decap_3 PHY_12167 ();
 sky130_fd_sc_hd__decap_3 PHY_12168 ();
 sky130_fd_sc_hd__decap_3 PHY_12169 ();
 sky130_fd_sc_hd__decap_3 PHY_12170 ();
 sky130_fd_sc_hd__decap_3 PHY_12171 ();
 sky130_fd_sc_hd__decap_3 PHY_12172 ();
 sky130_fd_sc_hd__decap_3 PHY_12173 ();
 sky130_fd_sc_hd__decap_3 PHY_12174 ();
 sky130_fd_sc_hd__decap_3 PHY_12175 ();
 sky130_fd_sc_hd__decap_3 PHY_12176 ();
 sky130_fd_sc_hd__decap_3 PHY_12177 ();
 sky130_fd_sc_hd__decap_3 PHY_12178 ();
 sky130_fd_sc_hd__decap_3 PHY_12179 ();
 sky130_fd_sc_hd__decap_3 PHY_12180 ();
 sky130_fd_sc_hd__decap_3 PHY_12181 ();
 sky130_fd_sc_hd__decap_3 PHY_12182 ();
 sky130_fd_sc_hd__decap_3 PHY_12183 ();
 sky130_fd_sc_hd__decap_3 PHY_12184 ();
 sky130_fd_sc_hd__decap_3 PHY_12185 ();
 sky130_fd_sc_hd__decap_3 PHY_12186 ();
 sky130_fd_sc_hd__decap_3 PHY_12187 ();
 sky130_fd_sc_hd__decap_3 PHY_12188 ();
 sky130_fd_sc_hd__decap_3 PHY_12189 ();
 sky130_fd_sc_hd__decap_3 PHY_12190 ();
 sky130_fd_sc_hd__decap_3 PHY_12191 ();
 sky130_fd_sc_hd__decap_3 PHY_12192 ();
 sky130_fd_sc_hd__decap_3 PHY_12193 ();
 sky130_fd_sc_hd__decap_3 PHY_12194 ();
 sky130_fd_sc_hd__decap_3 PHY_12195 ();
 sky130_fd_sc_hd__decap_3 PHY_12196 ();
 sky130_fd_sc_hd__decap_3 PHY_12197 ();
 sky130_fd_sc_hd__decap_3 PHY_12198 ();
 sky130_fd_sc_hd__decap_3 PHY_12199 ();
 sky130_fd_sc_hd__decap_3 PHY_12200 ();
 sky130_fd_sc_hd__decap_3 PHY_12201 ();
 sky130_fd_sc_hd__decap_3 PHY_12202 ();
 sky130_fd_sc_hd__decap_3 PHY_12203 ();
 sky130_fd_sc_hd__decap_3 PHY_12204 ();
 sky130_fd_sc_hd__decap_3 PHY_12205 ();
 sky130_fd_sc_hd__decap_3 PHY_12206 ();
 sky130_fd_sc_hd__decap_3 PHY_12207 ();
 sky130_fd_sc_hd__decap_3 PHY_12208 ();
 sky130_fd_sc_hd__decap_3 PHY_12209 ();
 sky130_fd_sc_hd__decap_3 PHY_12210 ();
 sky130_fd_sc_hd__decap_3 PHY_12211 ();
 sky130_fd_sc_hd__decap_3 PHY_12212 ();
 sky130_fd_sc_hd__decap_3 PHY_12213 ();
 sky130_fd_sc_hd__decap_3 PHY_12214 ();
 sky130_fd_sc_hd__decap_3 PHY_12215 ();
 sky130_fd_sc_hd__decap_3 PHY_12216 ();
 sky130_fd_sc_hd__decap_3 PHY_12217 ();
 sky130_fd_sc_hd__decap_3 PHY_12218 ();
 sky130_fd_sc_hd__decap_3 PHY_12219 ();
 sky130_fd_sc_hd__decap_3 PHY_12220 ();
 sky130_fd_sc_hd__decap_3 PHY_12221 ();
 sky130_fd_sc_hd__decap_3 PHY_12222 ();
 sky130_fd_sc_hd__decap_3 PHY_12223 ();
 sky130_fd_sc_hd__decap_3 PHY_12224 ();
 sky130_fd_sc_hd__decap_3 PHY_12225 ();
 sky130_fd_sc_hd__decap_3 PHY_12226 ();
 sky130_fd_sc_hd__decap_3 PHY_12227 ();
 sky130_fd_sc_hd__decap_3 PHY_12228 ();
 sky130_fd_sc_hd__decap_3 PHY_12229 ();
 sky130_fd_sc_hd__decap_3 PHY_12230 ();
 sky130_fd_sc_hd__decap_3 PHY_12231 ();
 sky130_fd_sc_hd__decap_3 PHY_12232 ();
 sky130_fd_sc_hd__decap_3 PHY_12233 ();
 sky130_fd_sc_hd__decap_3 PHY_12234 ();
 sky130_fd_sc_hd__decap_3 PHY_12235 ();
 sky130_fd_sc_hd__decap_3 PHY_12236 ();
 sky130_fd_sc_hd__decap_3 PHY_12237 ();
 sky130_fd_sc_hd__decap_3 PHY_12238 ();
 sky130_fd_sc_hd__decap_3 PHY_12239 ();
 sky130_fd_sc_hd__decap_3 PHY_12240 ();
 sky130_fd_sc_hd__decap_3 PHY_12241 ();
 sky130_fd_sc_hd__decap_3 PHY_12242 ();
 sky130_fd_sc_hd__decap_3 PHY_12243 ();
 sky130_fd_sc_hd__decap_3 PHY_12244 ();
 sky130_fd_sc_hd__decap_3 PHY_12245 ();
 sky130_fd_sc_hd__decap_3 PHY_12246 ();
 sky130_fd_sc_hd__decap_3 PHY_12247 ();
 sky130_fd_sc_hd__decap_3 PHY_12248 ();
 sky130_fd_sc_hd__decap_3 PHY_12249 ();
 sky130_fd_sc_hd__decap_3 PHY_12250 ();
 sky130_fd_sc_hd__decap_3 PHY_12251 ();
 sky130_fd_sc_hd__decap_3 PHY_12252 ();
 sky130_fd_sc_hd__decap_3 PHY_12253 ();
 sky130_fd_sc_hd__decap_3 PHY_12254 ();
 sky130_fd_sc_hd__decap_3 PHY_12255 ();
 sky130_fd_sc_hd__decap_3 PHY_12256 ();
 sky130_fd_sc_hd__decap_3 PHY_12257 ();
 sky130_fd_sc_hd__decap_3 PHY_12258 ();
 sky130_fd_sc_hd__decap_3 PHY_12259 ();
 sky130_fd_sc_hd__decap_3 PHY_12260 ();
 sky130_fd_sc_hd__decap_3 PHY_12261 ();
 sky130_fd_sc_hd__decap_3 PHY_12262 ();
 sky130_fd_sc_hd__decap_3 PHY_12263 ();
 sky130_fd_sc_hd__decap_3 PHY_12264 ();
 sky130_fd_sc_hd__decap_3 PHY_12265 ();
 sky130_fd_sc_hd__decap_3 PHY_12266 ();
 sky130_fd_sc_hd__decap_3 PHY_12267 ();
 sky130_fd_sc_hd__decap_3 PHY_12268 ();
 sky130_fd_sc_hd__decap_3 PHY_12269 ();
 sky130_fd_sc_hd__decap_3 PHY_12270 ();
 sky130_fd_sc_hd__decap_3 PHY_12271 ();
 sky130_fd_sc_hd__decap_3 PHY_12272 ();
 sky130_fd_sc_hd__decap_3 PHY_12273 ();
 sky130_fd_sc_hd__decap_3 PHY_12274 ();
 sky130_fd_sc_hd__decap_3 PHY_12275 ();
 sky130_fd_sc_hd__decap_3 PHY_12276 ();
 sky130_fd_sc_hd__decap_3 PHY_12277 ();
 sky130_fd_sc_hd__decap_3 PHY_12278 ();
 sky130_fd_sc_hd__decap_3 PHY_12279 ();
 sky130_fd_sc_hd__decap_3 PHY_12280 ();
 sky130_fd_sc_hd__decap_3 PHY_12281 ();
 sky130_fd_sc_hd__decap_3 PHY_12282 ();
 sky130_fd_sc_hd__decap_3 PHY_12283 ();
 sky130_fd_sc_hd__decap_3 PHY_12284 ();
 sky130_fd_sc_hd__decap_3 PHY_12285 ();
 sky130_fd_sc_hd__decap_3 PHY_12286 ();
 sky130_fd_sc_hd__decap_3 PHY_12287 ();
 sky130_fd_sc_hd__decap_3 PHY_12288 ();
 sky130_fd_sc_hd__decap_3 PHY_12289 ();
 sky130_fd_sc_hd__decap_3 PHY_12290 ();
 sky130_fd_sc_hd__decap_3 PHY_12291 ();
 sky130_fd_sc_hd__decap_3 PHY_12292 ();
 sky130_fd_sc_hd__decap_3 PHY_12293 ();
 sky130_fd_sc_hd__decap_3 PHY_12294 ();
 sky130_fd_sc_hd__decap_3 PHY_12295 ();
 sky130_fd_sc_hd__decap_3 PHY_12296 ();
 sky130_fd_sc_hd__decap_3 PHY_12297 ();
 sky130_fd_sc_hd__decap_3 PHY_12298 ();
 sky130_fd_sc_hd__decap_3 PHY_12299 ();
 sky130_fd_sc_hd__decap_3 PHY_12300 ();
 sky130_fd_sc_hd__decap_3 PHY_12301 ();
 sky130_fd_sc_hd__decap_3 PHY_12302 ();
 sky130_fd_sc_hd__decap_3 PHY_12303 ();
 sky130_fd_sc_hd__decap_3 PHY_12304 ();
 sky130_fd_sc_hd__decap_3 PHY_12305 ();
 sky130_fd_sc_hd__decap_3 PHY_12306 ();
 sky130_fd_sc_hd__decap_3 PHY_12307 ();
 sky130_fd_sc_hd__decap_3 PHY_12308 ();
 sky130_fd_sc_hd__decap_3 PHY_12309 ();
 sky130_fd_sc_hd__decap_3 PHY_12310 ();
 sky130_fd_sc_hd__decap_3 PHY_12311 ();
 sky130_fd_sc_hd__decap_3 PHY_12312 ();
 sky130_fd_sc_hd__decap_3 PHY_12313 ();
 sky130_fd_sc_hd__decap_3 PHY_12314 ();
 sky130_fd_sc_hd__decap_3 PHY_12315 ();
 sky130_fd_sc_hd__decap_3 PHY_12316 ();
 sky130_fd_sc_hd__decap_3 PHY_12317 ();
 sky130_fd_sc_hd__decap_3 PHY_12318 ();
 sky130_fd_sc_hd__decap_3 PHY_12319 ();
 sky130_fd_sc_hd__decap_3 PHY_12320 ();
 sky130_fd_sc_hd__decap_3 PHY_12321 ();
 sky130_fd_sc_hd__decap_3 PHY_12322 ();
 sky130_fd_sc_hd__decap_3 PHY_12323 ();
 sky130_fd_sc_hd__decap_3 PHY_12324 ();
 sky130_fd_sc_hd__decap_3 PHY_12325 ();
 sky130_fd_sc_hd__decap_3 PHY_12326 ();
 sky130_fd_sc_hd__decap_3 PHY_12327 ();
 sky130_fd_sc_hd__decap_3 PHY_12328 ();
 sky130_fd_sc_hd__decap_3 PHY_12329 ();
 sky130_fd_sc_hd__decap_3 PHY_12330 ();
 sky130_fd_sc_hd__decap_3 PHY_12331 ();
 sky130_fd_sc_hd__decap_3 PHY_12332 ();
 sky130_fd_sc_hd__decap_3 PHY_12333 ();
 sky130_fd_sc_hd__decap_3 PHY_12334 ();
 sky130_fd_sc_hd__decap_3 PHY_12335 ();
 sky130_fd_sc_hd__decap_3 PHY_12336 ();
 sky130_fd_sc_hd__decap_3 PHY_12337 ();
 sky130_fd_sc_hd__decap_3 PHY_12338 ();
 sky130_fd_sc_hd__decap_3 PHY_12339 ();
 sky130_fd_sc_hd__decap_3 PHY_12340 ();
 sky130_fd_sc_hd__decap_3 PHY_12341 ();
 sky130_fd_sc_hd__decap_3 PHY_12342 ();
 sky130_fd_sc_hd__decap_3 PHY_12343 ();
 sky130_fd_sc_hd__decap_3 PHY_12344 ();
 sky130_fd_sc_hd__decap_3 PHY_12345 ();
 sky130_fd_sc_hd__decap_3 PHY_12346 ();
 sky130_fd_sc_hd__decap_3 PHY_12347 ();
 sky130_fd_sc_hd__decap_3 PHY_12348 ();
 sky130_fd_sc_hd__decap_3 PHY_12349 ();
 sky130_fd_sc_hd__decap_3 PHY_12350 ();
 sky130_fd_sc_hd__decap_3 PHY_12351 ();
 sky130_fd_sc_hd__decap_3 PHY_12352 ();
 sky130_fd_sc_hd__decap_3 PHY_12353 ();
 sky130_fd_sc_hd__decap_3 PHY_12354 ();
 sky130_fd_sc_hd__decap_3 PHY_12355 ();
 sky130_fd_sc_hd__decap_3 PHY_12356 ();
 sky130_fd_sc_hd__decap_3 PHY_12357 ();
 sky130_fd_sc_hd__decap_3 PHY_12358 ();
 sky130_fd_sc_hd__decap_3 PHY_12359 ();
 sky130_fd_sc_hd__decap_3 PHY_12360 ();
 sky130_fd_sc_hd__decap_3 PHY_12361 ();
 sky130_fd_sc_hd__decap_3 PHY_12362 ();
 sky130_fd_sc_hd__decap_3 PHY_12363 ();
 sky130_fd_sc_hd__decap_3 PHY_12364 ();
 sky130_fd_sc_hd__decap_3 PHY_12365 ();
 sky130_fd_sc_hd__decap_3 PHY_12366 ();
 sky130_fd_sc_hd__decap_3 PHY_12367 ();
 sky130_fd_sc_hd__decap_3 PHY_12368 ();
 sky130_fd_sc_hd__decap_3 PHY_12369 ();
 sky130_fd_sc_hd__decap_3 PHY_12370 ();
 sky130_fd_sc_hd__decap_3 PHY_12371 ();
 sky130_fd_sc_hd__decap_3 PHY_12372 ();
 sky130_fd_sc_hd__decap_3 PHY_12373 ();
 sky130_fd_sc_hd__decap_3 PHY_12374 ();
 sky130_fd_sc_hd__decap_3 PHY_12375 ();
 sky130_fd_sc_hd__decap_3 PHY_12376 ();
 sky130_fd_sc_hd__decap_3 PHY_12377 ();
 sky130_fd_sc_hd__decap_3 PHY_12378 ();
 sky130_fd_sc_hd__decap_3 PHY_12379 ();
 sky130_fd_sc_hd__decap_3 PHY_12380 ();
 sky130_fd_sc_hd__decap_3 PHY_12381 ();
 sky130_fd_sc_hd__decap_3 PHY_12382 ();
 sky130_fd_sc_hd__decap_3 PHY_12383 ();
 sky130_fd_sc_hd__decap_3 PHY_12384 ();
 sky130_fd_sc_hd__decap_3 PHY_12385 ();
 sky130_fd_sc_hd__decap_3 PHY_12386 ();
 sky130_fd_sc_hd__decap_3 PHY_12387 ();
 sky130_fd_sc_hd__decap_3 PHY_12388 ();
 sky130_fd_sc_hd__decap_3 PHY_12389 ();
 sky130_fd_sc_hd__decap_3 PHY_12390 ();
 sky130_fd_sc_hd__decap_3 PHY_12391 ();
 sky130_fd_sc_hd__decap_3 PHY_12392 ();
 sky130_fd_sc_hd__decap_3 PHY_12393 ();
 sky130_fd_sc_hd__decap_3 PHY_12394 ();
 sky130_fd_sc_hd__decap_3 PHY_12395 ();
 sky130_fd_sc_hd__decap_3 PHY_12396 ();
 sky130_fd_sc_hd__decap_3 PHY_12397 ();
 sky130_fd_sc_hd__decap_3 PHY_12398 ();
 sky130_fd_sc_hd__decap_3 PHY_12399 ();
 sky130_fd_sc_hd__decap_3 PHY_12400 ();
 sky130_fd_sc_hd__decap_3 PHY_12401 ();
 sky130_fd_sc_hd__decap_3 PHY_12402 ();
 sky130_fd_sc_hd__decap_3 PHY_12403 ();
 sky130_fd_sc_hd__decap_3 PHY_12404 ();
 sky130_fd_sc_hd__decap_3 PHY_12405 ();
 sky130_fd_sc_hd__decap_3 PHY_12406 ();
 sky130_fd_sc_hd__decap_3 PHY_12407 ();
 sky130_fd_sc_hd__decap_3 PHY_12408 ();
 sky130_fd_sc_hd__decap_3 PHY_12409 ();
 sky130_fd_sc_hd__decap_3 PHY_12410 ();
 sky130_fd_sc_hd__decap_3 PHY_12411 ();
 sky130_fd_sc_hd__decap_3 PHY_12412 ();
 sky130_fd_sc_hd__decap_3 PHY_12413 ();
 sky130_fd_sc_hd__decap_3 PHY_12414 ();
 sky130_fd_sc_hd__decap_3 PHY_12415 ();
 sky130_fd_sc_hd__decap_3 PHY_12416 ();
 sky130_fd_sc_hd__decap_3 PHY_12417 ();
 sky130_fd_sc_hd__decap_3 PHY_12418 ();
 sky130_fd_sc_hd__decap_3 PHY_12419 ();
 sky130_fd_sc_hd__decap_3 PHY_12420 ();
 sky130_fd_sc_hd__decap_3 PHY_12421 ();
 sky130_fd_sc_hd__decap_3 PHY_12422 ();
 sky130_fd_sc_hd__decap_3 PHY_12423 ();
 sky130_fd_sc_hd__decap_3 PHY_12424 ();
 sky130_fd_sc_hd__decap_3 PHY_12425 ();
 sky130_fd_sc_hd__decap_3 PHY_12426 ();
 sky130_fd_sc_hd__decap_3 PHY_12427 ();
 sky130_fd_sc_hd__decap_3 PHY_12428 ();
 sky130_fd_sc_hd__decap_3 PHY_12429 ();
 sky130_fd_sc_hd__decap_3 PHY_12430 ();
 sky130_fd_sc_hd__decap_3 PHY_12431 ();
 sky130_fd_sc_hd__decap_3 PHY_12432 ();
 sky130_fd_sc_hd__decap_3 PHY_12433 ();
 sky130_fd_sc_hd__decap_3 PHY_12434 ();
 sky130_fd_sc_hd__decap_3 PHY_12435 ();
 sky130_fd_sc_hd__decap_3 PHY_12436 ();
 sky130_fd_sc_hd__decap_3 PHY_12437 ();
 sky130_fd_sc_hd__decap_3 PHY_12438 ();
 sky130_fd_sc_hd__decap_3 PHY_12439 ();
 sky130_fd_sc_hd__decap_3 PHY_12440 ();
 sky130_fd_sc_hd__decap_3 PHY_12441 ();
 sky130_fd_sc_hd__decap_3 PHY_12442 ();
 sky130_fd_sc_hd__decap_3 PHY_12443 ();
 sky130_fd_sc_hd__decap_3 PHY_12444 ();
 sky130_fd_sc_hd__decap_3 PHY_12445 ();
 sky130_fd_sc_hd__decap_3 PHY_12446 ();
 sky130_fd_sc_hd__decap_3 PHY_12447 ();
 sky130_fd_sc_hd__decap_3 PHY_12448 ();
 sky130_fd_sc_hd__decap_3 PHY_12449 ();
 sky130_fd_sc_hd__decap_3 PHY_12450 ();
 sky130_fd_sc_hd__decap_3 PHY_12451 ();
 sky130_fd_sc_hd__decap_3 PHY_12452 ();
 sky130_fd_sc_hd__decap_3 PHY_12453 ();
 sky130_fd_sc_hd__decap_3 PHY_12454 ();
 sky130_fd_sc_hd__decap_3 PHY_12455 ();
 sky130_fd_sc_hd__decap_3 PHY_12456 ();
 sky130_fd_sc_hd__decap_3 PHY_12457 ();
 sky130_fd_sc_hd__decap_3 PHY_12458 ();
 sky130_fd_sc_hd__decap_3 PHY_12459 ();
 sky130_fd_sc_hd__decap_3 PHY_12460 ();
 sky130_fd_sc_hd__decap_3 PHY_12461 ();
 sky130_fd_sc_hd__decap_3 PHY_12462 ();
 sky130_fd_sc_hd__decap_3 PHY_12463 ();
 sky130_fd_sc_hd__decap_3 PHY_12464 ();
 sky130_fd_sc_hd__decap_3 PHY_12465 ();
 sky130_fd_sc_hd__decap_3 PHY_12466 ();
 sky130_fd_sc_hd__decap_3 PHY_12467 ();
 sky130_fd_sc_hd__decap_3 PHY_12468 ();
 sky130_fd_sc_hd__decap_3 PHY_12469 ();
 sky130_fd_sc_hd__decap_3 PHY_12470 ();
 sky130_fd_sc_hd__decap_3 PHY_12471 ();
 sky130_fd_sc_hd__decap_3 PHY_12472 ();
 sky130_fd_sc_hd__decap_3 PHY_12473 ();
 sky130_fd_sc_hd__decap_3 PHY_12474 ();
 sky130_fd_sc_hd__decap_3 PHY_12475 ();
 sky130_fd_sc_hd__decap_3 PHY_12476 ();
 sky130_fd_sc_hd__decap_3 PHY_12477 ();
 sky130_fd_sc_hd__decap_3 PHY_12478 ();
 sky130_fd_sc_hd__decap_3 PHY_12479 ();
 sky130_fd_sc_hd__decap_3 PHY_12480 ();
 sky130_fd_sc_hd__decap_3 PHY_12481 ();
 sky130_fd_sc_hd__decap_3 PHY_12482 ();
 sky130_fd_sc_hd__decap_3 PHY_12483 ();
 sky130_fd_sc_hd__decap_3 PHY_12484 ();
 sky130_fd_sc_hd__decap_3 PHY_12485 ();
 sky130_fd_sc_hd__decap_3 PHY_12486 ();
 sky130_fd_sc_hd__decap_3 PHY_12487 ();
 sky130_fd_sc_hd__decap_3 PHY_12488 ();
 sky130_fd_sc_hd__decap_3 PHY_12489 ();
 sky130_fd_sc_hd__decap_3 PHY_12490 ();
 sky130_fd_sc_hd__decap_3 PHY_12491 ();
 sky130_fd_sc_hd__decap_3 PHY_12492 ();
 sky130_fd_sc_hd__decap_3 PHY_12493 ();
 sky130_fd_sc_hd__decap_3 PHY_12494 ();
 sky130_fd_sc_hd__decap_3 PHY_12495 ();
 sky130_fd_sc_hd__decap_3 PHY_12496 ();
 sky130_fd_sc_hd__decap_3 PHY_12497 ();
 sky130_fd_sc_hd__decap_3 PHY_12498 ();
 sky130_fd_sc_hd__decap_3 PHY_12499 ();
 sky130_fd_sc_hd__decap_3 PHY_12500 ();
 sky130_fd_sc_hd__decap_3 PHY_12501 ();
 sky130_fd_sc_hd__decap_3 PHY_12502 ();
 sky130_fd_sc_hd__decap_3 PHY_12503 ();
 sky130_fd_sc_hd__decap_3 PHY_12504 ();
 sky130_fd_sc_hd__decap_3 PHY_12505 ();
 sky130_fd_sc_hd__decap_3 PHY_12506 ();
 sky130_fd_sc_hd__decap_3 PHY_12507 ();
 sky130_fd_sc_hd__decap_3 PHY_12508 ();
 sky130_fd_sc_hd__decap_3 PHY_12509 ();
 sky130_fd_sc_hd__decap_3 PHY_12510 ();
 sky130_fd_sc_hd__decap_3 PHY_12511 ();
 sky130_fd_sc_hd__decap_3 PHY_12512 ();
 sky130_fd_sc_hd__decap_3 PHY_12513 ();
 sky130_fd_sc_hd__decap_3 PHY_12514 ();
 sky130_fd_sc_hd__decap_3 PHY_12515 ();
 sky130_fd_sc_hd__decap_3 PHY_12516 ();
 sky130_fd_sc_hd__decap_3 PHY_12517 ();
 sky130_fd_sc_hd__decap_3 PHY_12518 ();
 sky130_fd_sc_hd__decap_3 PHY_12519 ();
 sky130_fd_sc_hd__decap_3 PHY_12520 ();
 sky130_fd_sc_hd__decap_3 PHY_12521 ();
 sky130_fd_sc_hd__decap_3 PHY_12522 ();
 sky130_fd_sc_hd__decap_3 PHY_12523 ();
 sky130_fd_sc_hd__decap_3 PHY_12524 ();
 sky130_fd_sc_hd__decap_3 PHY_12525 ();
 sky130_fd_sc_hd__decap_3 PHY_12526 ();
 sky130_fd_sc_hd__decap_3 PHY_12527 ();
 sky130_fd_sc_hd__decap_3 PHY_12528 ();
 sky130_fd_sc_hd__decap_3 PHY_12529 ();
 sky130_fd_sc_hd__decap_3 PHY_12530 ();
 sky130_fd_sc_hd__decap_3 PHY_12531 ();
 sky130_fd_sc_hd__decap_3 PHY_12532 ();
 sky130_fd_sc_hd__decap_3 PHY_12533 ();
 sky130_fd_sc_hd__decap_3 PHY_12534 ();
 sky130_fd_sc_hd__decap_3 PHY_12535 ();
 sky130_fd_sc_hd__decap_3 PHY_12536 ();
 sky130_fd_sc_hd__decap_3 PHY_12537 ();
 sky130_fd_sc_hd__decap_3 PHY_12538 ();
 sky130_fd_sc_hd__decap_3 PHY_12539 ();
 sky130_fd_sc_hd__decap_3 PHY_12540 ();
 sky130_fd_sc_hd__decap_3 PHY_12541 ();
 sky130_fd_sc_hd__decap_3 PHY_12542 ();
 sky130_fd_sc_hd__decap_3 PHY_12543 ();
 sky130_fd_sc_hd__decap_3 PHY_12544 ();
 sky130_fd_sc_hd__decap_3 PHY_12545 ();
 sky130_fd_sc_hd__decap_3 PHY_12546 ();
 sky130_fd_sc_hd__decap_3 PHY_12547 ();
 sky130_fd_sc_hd__decap_3 PHY_12548 ();
 sky130_fd_sc_hd__decap_3 PHY_12549 ();
 sky130_fd_sc_hd__decap_3 PHY_12550 ();
 sky130_fd_sc_hd__decap_3 PHY_12551 ();
 sky130_fd_sc_hd__decap_3 PHY_12552 ();
 sky130_fd_sc_hd__decap_3 PHY_12553 ();
 sky130_fd_sc_hd__decap_3 PHY_12554 ();
 sky130_fd_sc_hd__decap_3 PHY_12555 ();
 sky130_fd_sc_hd__decap_3 PHY_12556 ();
 sky130_fd_sc_hd__decap_3 PHY_12557 ();
 sky130_fd_sc_hd__decap_3 PHY_12558 ();
 sky130_fd_sc_hd__decap_3 PHY_12559 ();
 sky130_fd_sc_hd__decap_3 PHY_12560 ();
 sky130_fd_sc_hd__decap_3 PHY_12561 ();
 sky130_fd_sc_hd__decap_3 PHY_12562 ();
 sky130_fd_sc_hd__decap_3 PHY_12563 ();
 sky130_fd_sc_hd__decap_3 PHY_12564 ();
 sky130_fd_sc_hd__decap_3 PHY_12565 ();
 sky130_fd_sc_hd__decap_3 PHY_12566 ();
 sky130_fd_sc_hd__decap_3 PHY_12567 ();
 sky130_fd_sc_hd__decap_3 PHY_12568 ();
 sky130_fd_sc_hd__decap_3 PHY_12569 ();
 sky130_fd_sc_hd__decap_3 PHY_12570 ();
 sky130_fd_sc_hd__decap_3 PHY_12571 ();
 sky130_fd_sc_hd__decap_3 PHY_12572 ();
 sky130_fd_sc_hd__decap_3 PHY_12573 ();
 sky130_fd_sc_hd__decap_3 PHY_12574 ();
 sky130_fd_sc_hd__decap_3 PHY_12575 ();
 sky130_fd_sc_hd__decap_3 PHY_12576 ();
 sky130_fd_sc_hd__decap_3 PHY_12577 ();
 sky130_fd_sc_hd__decap_3 PHY_12578 ();
 sky130_fd_sc_hd__decap_3 PHY_12579 ();
 sky130_fd_sc_hd__decap_3 PHY_12580 ();
 sky130_fd_sc_hd__decap_3 PHY_12581 ();
 sky130_fd_sc_hd__decap_3 PHY_12582 ();
 sky130_fd_sc_hd__decap_3 PHY_12583 ();
 sky130_fd_sc_hd__decap_3 PHY_12584 ();
 sky130_fd_sc_hd__decap_3 PHY_12585 ();
 sky130_fd_sc_hd__decap_3 PHY_12586 ();
 sky130_fd_sc_hd__decap_3 PHY_12587 ();
 sky130_fd_sc_hd__decap_3 PHY_12588 ();
 sky130_fd_sc_hd__decap_3 PHY_12589 ();
 sky130_fd_sc_hd__decap_3 PHY_12590 ();
 sky130_fd_sc_hd__decap_3 PHY_12591 ();
 sky130_fd_sc_hd__decap_3 PHY_12592 ();
 sky130_fd_sc_hd__decap_3 PHY_12593 ();
 sky130_fd_sc_hd__decap_3 PHY_12594 ();
 sky130_fd_sc_hd__decap_3 PHY_12595 ();
 sky130_fd_sc_hd__decap_3 PHY_12596 ();
 sky130_fd_sc_hd__decap_3 PHY_12597 ();
 sky130_fd_sc_hd__decap_3 PHY_12598 ();
 sky130_fd_sc_hd__decap_3 PHY_12599 ();
 sky130_fd_sc_hd__decap_3 PHY_12600 ();
 sky130_fd_sc_hd__decap_3 PHY_12601 ();
 sky130_fd_sc_hd__decap_3 PHY_12602 ();
 sky130_fd_sc_hd__decap_3 PHY_12603 ();
 sky130_fd_sc_hd__decap_3 PHY_12604 ();
 sky130_fd_sc_hd__decap_3 PHY_12605 ();
 sky130_fd_sc_hd__decap_3 PHY_12606 ();
 sky130_fd_sc_hd__decap_3 PHY_12607 ();
 sky130_fd_sc_hd__decap_3 PHY_12608 ();
 sky130_fd_sc_hd__decap_3 PHY_12609 ();
 sky130_fd_sc_hd__decap_3 PHY_12610 ();
 sky130_fd_sc_hd__decap_3 PHY_12611 ();
 sky130_fd_sc_hd__decap_3 PHY_12612 ();
 sky130_fd_sc_hd__decap_3 PHY_12613 ();
 sky130_fd_sc_hd__decap_3 PHY_12614 ();
 sky130_fd_sc_hd__decap_3 PHY_12615 ();
 sky130_fd_sc_hd__decap_3 PHY_12616 ();
 sky130_fd_sc_hd__decap_3 PHY_12617 ();
 sky130_fd_sc_hd__decap_3 PHY_12618 ();
 sky130_fd_sc_hd__decap_3 PHY_12619 ();
 sky130_fd_sc_hd__decap_3 PHY_12620 ();
 sky130_fd_sc_hd__decap_3 PHY_12621 ();
 sky130_fd_sc_hd__decap_3 PHY_12622 ();
 sky130_fd_sc_hd__decap_3 PHY_12623 ();
 sky130_fd_sc_hd__decap_3 PHY_12624 ();
 sky130_fd_sc_hd__decap_3 PHY_12625 ();
 sky130_fd_sc_hd__decap_3 PHY_12626 ();
 sky130_fd_sc_hd__decap_3 PHY_12627 ();
 sky130_fd_sc_hd__decap_3 PHY_12628 ();
 sky130_fd_sc_hd__decap_3 PHY_12629 ();
 sky130_fd_sc_hd__decap_3 PHY_12630 ();
 sky130_fd_sc_hd__decap_3 PHY_12631 ();
 sky130_fd_sc_hd__decap_3 PHY_12632 ();
 sky130_fd_sc_hd__decap_3 PHY_12633 ();
 sky130_fd_sc_hd__decap_3 PHY_12634 ();
 sky130_fd_sc_hd__decap_3 PHY_12635 ();
 sky130_fd_sc_hd__decap_3 PHY_12636 ();
 sky130_fd_sc_hd__decap_3 PHY_12637 ();
 sky130_fd_sc_hd__decap_3 PHY_12638 ();
 sky130_fd_sc_hd__decap_3 PHY_12639 ();
 sky130_fd_sc_hd__decap_3 PHY_12640 ();
 sky130_fd_sc_hd__decap_3 PHY_12641 ();
 sky130_fd_sc_hd__decap_3 PHY_12642 ();
 sky130_fd_sc_hd__decap_3 PHY_12643 ();
 sky130_fd_sc_hd__decap_3 PHY_12644 ();
 sky130_fd_sc_hd__decap_3 PHY_12645 ();
 sky130_fd_sc_hd__decap_3 PHY_12646 ();
 sky130_fd_sc_hd__decap_3 PHY_12647 ();
 sky130_fd_sc_hd__decap_3 PHY_12648 ();
 sky130_fd_sc_hd__decap_3 PHY_12649 ();
 sky130_fd_sc_hd__decap_3 PHY_12650 ();
 sky130_fd_sc_hd__decap_3 PHY_12651 ();
 sky130_fd_sc_hd__decap_3 PHY_12652 ();
 sky130_fd_sc_hd__decap_3 PHY_12653 ();
 sky130_fd_sc_hd__decap_3 PHY_12654 ();
 sky130_fd_sc_hd__decap_3 PHY_12655 ();
 sky130_fd_sc_hd__decap_3 PHY_12656 ();
 sky130_fd_sc_hd__decap_3 PHY_12657 ();
 sky130_fd_sc_hd__decap_3 PHY_12658 ();
 sky130_fd_sc_hd__decap_3 PHY_12659 ();
 sky130_fd_sc_hd__decap_3 PHY_12660 ();
 sky130_fd_sc_hd__decap_3 PHY_12661 ();
 sky130_fd_sc_hd__decap_3 PHY_12662 ();
 sky130_fd_sc_hd__decap_3 PHY_12663 ();
 sky130_fd_sc_hd__decap_3 PHY_12664 ();
 sky130_fd_sc_hd__decap_3 PHY_12665 ();
 sky130_fd_sc_hd__decap_3 PHY_12666 ();
 sky130_fd_sc_hd__decap_3 PHY_12667 ();
 sky130_fd_sc_hd__decap_3 PHY_12668 ();
 sky130_fd_sc_hd__decap_3 PHY_12669 ();
 sky130_fd_sc_hd__decap_3 PHY_12670 ();
 sky130_fd_sc_hd__decap_3 PHY_12671 ();
 sky130_fd_sc_hd__decap_3 PHY_12672 ();
 sky130_fd_sc_hd__decap_3 PHY_12673 ();
 sky130_fd_sc_hd__decap_3 PHY_12674 ();
 sky130_fd_sc_hd__decap_3 PHY_12675 ();
 sky130_fd_sc_hd__decap_3 PHY_12676 ();
 sky130_fd_sc_hd__decap_3 PHY_12677 ();
 sky130_fd_sc_hd__decap_3 PHY_12678 ();
 sky130_fd_sc_hd__decap_3 PHY_12679 ();
 sky130_fd_sc_hd__decap_3 PHY_12680 ();
 sky130_fd_sc_hd__decap_3 PHY_12681 ();
 sky130_fd_sc_hd__decap_3 PHY_12682 ();
 sky130_fd_sc_hd__decap_3 PHY_12683 ();
 sky130_fd_sc_hd__decap_3 PHY_12684 ();
 sky130_fd_sc_hd__decap_3 PHY_12685 ();
 sky130_fd_sc_hd__decap_3 PHY_12686 ();
 sky130_fd_sc_hd__decap_3 PHY_12687 ();
 sky130_fd_sc_hd__decap_3 PHY_12688 ();
 sky130_fd_sc_hd__decap_3 PHY_12689 ();
 sky130_fd_sc_hd__decap_3 PHY_12690 ();
 sky130_fd_sc_hd__decap_3 PHY_12691 ();
 sky130_fd_sc_hd__decap_3 PHY_12692 ();
 sky130_fd_sc_hd__decap_3 PHY_12693 ();
 sky130_fd_sc_hd__decap_3 PHY_12694 ();
 sky130_fd_sc_hd__decap_3 PHY_12695 ();
 sky130_fd_sc_hd__decap_3 PHY_12696 ();
 sky130_fd_sc_hd__decap_3 PHY_12697 ();
 sky130_fd_sc_hd__decap_3 PHY_12698 ();
 sky130_fd_sc_hd__decap_3 PHY_12699 ();
 sky130_fd_sc_hd__decap_3 PHY_12700 ();
 sky130_fd_sc_hd__decap_3 PHY_12701 ();
 sky130_fd_sc_hd__decap_3 PHY_12702 ();
 sky130_fd_sc_hd__decap_3 PHY_12703 ();
 sky130_fd_sc_hd__decap_3 PHY_12704 ();
 sky130_fd_sc_hd__decap_3 PHY_12705 ();
 sky130_fd_sc_hd__decap_3 PHY_12706 ();
 sky130_fd_sc_hd__decap_3 PHY_12707 ();
 sky130_fd_sc_hd__decap_3 PHY_12708 ();
 sky130_fd_sc_hd__decap_3 PHY_12709 ();
 sky130_fd_sc_hd__decap_3 PHY_12710 ();
 sky130_fd_sc_hd__decap_3 PHY_12711 ();
 sky130_fd_sc_hd__decap_3 PHY_12712 ();
 sky130_fd_sc_hd__decap_3 PHY_12713 ();
 sky130_fd_sc_hd__decap_3 PHY_12714 ();
 sky130_fd_sc_hd__decap_3 PHY_12715 ();
 sky130_fd_sc_hd__decap_3 PHY_12716 ();
 sky130_fd_sc_hd__decap_3 PHY_12717 ();
 sky130_fd_sc_hd__decap_3 PHY_12718 ();
 sky130_fd_sc_hd__decap_3 PHY_12719 ();
 sky130_fd_sc_hd__decap_3 PHY_12720 ();
 sky130_fd_sc_hd__decap_3 PHY_12721 ();
 sky130_fd_sc_hd__decap_3 PHY_12722 ();
 sky130_fd_sc_hd__decap_3 PHY_12723 ();
 sky130_fd_sc_hd__decap_3 PHY_12724 ();
 sky130_fd_sc_hd__decap_3 PHY_12725 ();
 sky130_fd_sc_hd__decap_3 PHY_12726 ();
 sky130_fd_sc_hd__decap_3 PHY_12727 ();
 sky130_fd_sc_hd__decap_3 PHY_12728 ();
 sky130_fd_sc_hd__decap_3 PHY_12729 ();
 sky130_fd_sc_hd__decap_3 PHY_12730 ();
 sky130_fd_sc_hd__decap_3 PHY_12731 ();
 sky130_fd_sc_hd__decap_3 PHY_12732 ();
 sky130_fd_sc_hd__decap_3 PHY_12733 ();
 sky130_fd_sc_hd__decap_3 PHY_12734 ();
 sky130_fd_sc_hd__decap_3 PHY_12735 ();
 sky130_fd_sc_hd__decap_3 PHY_12736 ();
 sky130_fd_sc_hd__decap_3 PHY_12737 ();
 sky130_fd_sc_hd__decap_3 PHY_12738 ();
 sky130_fd_sc_hd__decap_3 PHY_12739 ();
 sky130_fd_sc_hd__decap_3 PHY_12740 ();
 sky130_fd_sc_hd__decap_3 PHY_12741 ();
 sky130_fd_sc_hd__decap_3 PHY_12742 ();
 sky130_fd_sc_hd__decap_3 PHY_12743 ();
 sky130_fd_sc_hd__decap_3 PHY_12744 ();
 sky130_fd_sc_hd__decap_3 PHY_12745 ();
 sky130_fd_sc_hd__decap_3 PHY_12746 ();
 sky130_fd_sc_hd__decap_3 PHY_12747 ();
 sky130_fd_sc_hd__decap_3 PHY_12748 ();
 sky130_fd_sc_hd__decap_3 PHY_12749 ();
 sky130_fd_sc_hd__decap_3 PHY_12750 ();
 sky130_fd_sc_hd__decap_3 PHY_12751 ();
 sky130_fd_sc_hd__decap_3 PHY_12752 ();
 sky130_fd_sc_hd__decap_3 PHY_12753 ();
 sky130_fd_sc_hd__decap_3 PHY_12754 ();
 sky130_fd_sc_hd__decap_3 PHY_12755 ();
 sky130_fd_sc_hd__decap_3 PHY_12756 ();
 sky130_fd_sc_hd__decap_3 PHY_12757 ();
 sky130_fd_sc_hd__decap_3 PHY_12758 ();
 sky130_fd_sc_hd__decap_3 PHY_12759 ();
 sky130_fd_sc_hd__decap_3 PHY_12760 ();
 sky130_fd_sc_hd__decap_3 PHY_12761 ();
 sky130_fd_sc_hd__decap_3 PHY_12762 ();
 sky130_fd_sc_hd__decap_3 PHY_12763 ();
 sky130_fd_sc_hd__decap_3 PHY_12764 ();
 sky130_fd_sc_hd__decap_3 PHY_12765 ();
 sky130_fd_sc_hd__decap_3 PHY_12766 ();
 sky130_fd_sc_hd__decap_3 PHY_12767 ();
 sky130_fd_sc_hd__decap_3 PHY_12768 ();
 sky130_fd_sc_hd__decap_3 PHY_12769 ();
 sky130_fd_sc_hd__decap_3 PHY_12770 ();
 sky130_fd_sc_hd__decap_3 PHY_12771 ();
 sky130_fd_sc_hd__decap_3 PHY_12772 ();
 sky130_fd_sc_hd__decap_3 PHY_12773 ();
 sky130_fd_sc_hd__decap_3 PHY_12774 ();
 sky130_fd_sc_hd__decap_3 PHY_12775 ();
 sky130_fd_sc_hd__decap_3 PHY_12776 ();
 sky130_fd_sc_hd__decap_3 PHY_12777 ();
 sky130_fd_sc_hd__decap_3 PHY_12778 ();
 sky130_fd_sc_hd__decap_3 PHY_12779 ();
 sky130_fd_sc_hd__decap_3 PHY_12780 ();
 sky130_fd_sc_hd__decap_3 PHY_12781 ();
 sky130_fd_sc_hd__decap_3 PHY_12782 ();
 sky130_fd_sc_hd__decap_3 PHY_12783 ();
 sky130_fd_sc_hd__decap_3 PHY_12784 ();
 sky130_fd_sc_hd__decap_3 PHY_12785 ();
 sky130_fd_sc_hd__decap_3 PHY_12786 ();
 sky130_fd_sc_hd__decap_3 PHY_12787 ();
 sky130_fd_sc_hd__decap_3 PHY_12788 ();
 sky130_fd_sc_hd__decap_3 PHY_12789 ();
 sky130_fd_sc_hd__decap_3 PHY_12790 ();
 sky130_fd_sc_hd__decap_3 PHY_12791 ();
 sky130_fd_sc_hd__decap_3 PHY_12792 ();
 sky130_fd_sc_hd__decap_3 PHY_12793 ();
 sky130_fd_sc_hd__decap_3 PHY_12794 ();
 sky130_fd_sc_hd__decap_3 PHY_12795 ();
 sky130_fd_sc_hd__decap_3 PHY_12796 ();
 sky130_fd_sc_hd__decap_3 PHY_12797 ();
 sky130_fd_sc_hd__decap_3 PHY_12798 ();
 sky130_fd_sc_hd__decap_3 PHY_12799 ();
 sky130_fd_sc_hd__decap_3 PHY_12800 ();
 sky130_fd_sc_hd__decap_3 PHY_12801 ();
 sky130_fd_sc_hd__decap_3 PHY_12802 ();
 sky130_fd_sc_hd__decap_3 PHY_12803 ();
 sky130_fd_sc_hd__decap_3 PHY_12804 ();
 sky130_fd_sc_hd__decap_3 PHY_12805 ();
 sky130_fd_sc_hd__decap_3 PHY_12806 ();
 sky130_fd_sc_hd__decap_3 PHY_12807 ();
 sky130_fd_sc_hd__decap_3 PHY_12808 ();
 sky130_fd_sc_hd__decap_3 PHY_12809 ();
 sky130_fd_sc_hd__decap_3 PHY_12810 ();
 sky130_fd_sc_hd__decap_3 PHY_12811 ();
 sky130_fd_sc_hd__decap_3 PHY_12812 ();
 sky130_fd_sc_hd__decap_3 PHY_12813 ();
 sky130_fd_sc_hd__decap_3 PHY_12814 ();
 sky130_fd_sc_hd__decap_3 PHY_12815 ();
 sky130_fd_sc_hd__decap_3 PHY_12816 ();
 sky130_fd_sc_hd__decap_3 PHY_12817 ();
 sky130_fd_sc_hd__decap_3 PHY_12818 ();
 sky130_fd_sc_hd__decap_3 PHY_12819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23445 ();
 sky130_fd_sc_hd__buf_8 input1 (.A(inp_data[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input2 (.A(inp_data[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(inp_data[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input4 (.A(inp_data[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(inp_data[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input6 (.A(inp_data[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(inp_data[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input8 (.A(inp_data[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input9 (.A(inp_data[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(inp_data[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input11 (.A(inp_data[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(inp_data[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(inp_data[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input14 (.A(inp_data[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(inp_data[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_12 input16 (.A(inp_data[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(inp_load),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(inp_y_addr[0]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_16 input19 (.A(inp_y_addr[1]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(inp_y_addr[2]),
    .X(net20));
 sky130_fd_sc_hd__buf_6 input21 (.A(inp_y_addr[3]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_16 input22 (.A(out_load),
    .X(net22));
 sky130_fd_sc_hd__buf_12 input23 (.A(out_shift),
    .X(net23));
 sky130_fd_sc_hd__buf_12 input24 (.A(net327),
    .X(net24));
 sky130_fd_sc_hd__buf_12 input25 (.A(run),
    .X(net25));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(out_data[0]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(out_data[10]));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net28),
    .X(out_data[11]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(out_data[12]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(out_data[13]));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net31),
    .X(out_data[14]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(out_data[15]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(out_data[1]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(out_data[2]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(out_data[3]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(out_data[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(out_data[5]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(out_data[6]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(out_data[7]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(out_data[8]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(out_data[9]));
 sky130_fd_sc_hd__buf_2 wire42 (.A(net48),
    .X(net42));
 sky130_fd_sc_hd__buf_2 wire43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_2 max_cap44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_2 wire45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_2 wire46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_2 wire47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__buf_2 wire48 (.A(_01_),
    .X(net48));
 sky130_fd_sc_hd__buf_8 wire49 (.A(\cell_outs[6] ),
    .X(net49));
 sky130_fd_sc_hd__buf_12 wire50 (.A(net9),
    .X(net50));
 sky130_fd_sc_hd__buf_12 wire51 (.A(net7),
    .X(net51));
 sky130_fd_sc_hd__buf_12 load_slew52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_12 load_slew53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_12 load_slew54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_12 load_slew55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_12 load_slew56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__buf_12 load_slew57 (.A(net66),
    .X(net57));
 sky130_fd_sc_hd__buf_12 load_slew58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_12 load_slew59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_12 load_slew60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_12 load_slew61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__buf_12 load_slew62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_12 load_slew63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_12 load_slew64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_12 load_slew65 (.A(net25),
    .X(net65));
 sky130_fd_sc_hd__buf_12 load_slew66 (.A(net25),
    .X(net66));
 sky130_fd_sc_hd__buf_12 load_slew67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_12 load_slew68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_12 load_slew69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_12 load_slew70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_12 load_slew71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_12 load_slew72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_12 load_slew73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__buf_12 load_slew74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_12 load_slew75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_12 load_slew76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_12 load_slew77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_12 load_slew78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_12 load_slew79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_12 load_slew80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_12 load_slew81 (.A(net24),
    .X(net81));
 sky130_fd_sc_hd__buf_12 load_slew82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_12 load_slew83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_12 load_slew84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_12 load_slew85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_12 load_slew86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_12 load_slew87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_12 load_slew88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_12 load_slew89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_12 load_slew90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_12 load_slew91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_12 load_slew92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_12 load_slew93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_12 load_slew94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_12 load_slew95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_12 load_slew96 (.A(net23),
    .X(net96));
 sky130_fd_sc_hd__buf_12 load_slew97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_16 load_slew98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_16 load_slew99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 load_slew100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_16 load_slew101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_16 load_slew102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_16 load_slew103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_16 load_slew104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_16 load_slew105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_16 load_slew106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_16 load_slew107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_16 load_slew108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_16 load_slew109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_16 load_slew110 (.A(net115),
    .X(net110));
 sky130_fd_sc_hd__buf_12 load_slew111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_12 load_slew112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_12 load_slew113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_12 load_slew114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_12 load_slew115 (.A(net22),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(net20),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout117 (.A(net20),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net19),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(net19),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net18),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout121 (.A(net18),
    .X(net121));
 sky130_fd_sc_hd__buf_12 wire122 (.A(net1),
    .X(net122));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y0_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y0_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y0_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y0_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y0_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y1_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y1_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y1_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y10_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y10_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y10_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y11_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y11_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y11_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y12_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y12_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y12_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y13_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y13_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y13_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y14_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y14_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y14_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y15_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y15_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y15_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y15_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y15_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y15_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y2_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y2_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y2_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y3_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y3_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y3_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y4_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y4_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y4_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y5_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y5_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y5_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y6_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y6_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y6_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y7_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y7_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y7_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y8_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y8_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y8_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y9_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y9_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 arr_cell_x0_y9_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y0_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y0_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y0_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y15_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y15_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y15_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 arr_cell_x10_y15_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y0_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y0_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y0_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y15_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y15_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y15_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 arr_cell_x11_y15_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y0_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y0_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y0_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y15_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y15_194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y15_195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 arr_cell_x12_y15_196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y0_197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y0_198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y0_199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y15_200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y15_201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y15_202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 arr_cell_x13_y15_203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y0_204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y0_205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y0_206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y15_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y15_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y15_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 arr_cell_x14_y15_210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y0_211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y0_212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y0_213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y0_214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y0_215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y1_216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y1_217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y1_218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y10_219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y10_220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y10_221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y11_222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y11_223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y11_224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y12_225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y12_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y12_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y13_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y13_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y13_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y14_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y14_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y14_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y15_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y15_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y15_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y15_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y15_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y15_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y2_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y2_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y2_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y3_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y3_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y3_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y4_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y4_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y4_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y5_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y5_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y5_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y6_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y6_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y6_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y7_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y7_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y7_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y8_258 (.LO(net258));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y8_259 (.LO(net259));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y8_260 (.LO(net260));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y9_261 (.LO(net261));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y9_262 (.LO(net262));
 sky130_fd_sc_hd__conb_1 arr_cell_x15_y9_263 (.LO(net263));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y0_264 (.LO(net264));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y0_265 (.LO(net265));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y0_266 (.LO(net266));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y15_267 (.LO(net267));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y15_268 (.LO(net268));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y15_269 (.LO(net269));
 sky130_fd_sc_hd__conb_1 arr_cell_x1_y15_270 (.LO(net270));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y0_271 (.LO(net271));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y0_272 (.LO(net272));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y0_273 (.LO(net273));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y15_274 (.LO(net274));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y15_275 (.LO(net275));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y15_276 (.LO(net276));
 sky130_fd_sc_hd__conb_1 arr_cell_x2_y15_277 (.LO(net277));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y0_278 (.LO(net278));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y0_279 (.LO(net279));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y0_280 (.LO(net280));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y15_281 (.LO(net281));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y15_282 (.LO(net282));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y15_283 (.LO(net283));
 sky130_fd_sc_hd__conb_1 arr_cell_x3_y15_284 (.LO(net284));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y0_285 (.LO(net285));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y0_286 (.LO(net286));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y0_287 (.LO(net287));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y15_288 (.LO(net288));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y15_289 (.LO(net289));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y15_290 (.LO(net290));
 sky130_fd_sc_hd__conb_1 arr_cell_x4_y15_291 (.LO(net291));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y0_292 (.LO(net292));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y0_293 (.LO(net293));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y0_294 (.LO(net294));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y15_295 (.LO(net295));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y15_296 (.LO(net296));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y15_297 (.LO(net297));
 sky130_fd_sc_hd__conb_1 arr_cell_x5_y15_298 (.LO(net298));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y0_299 (.LO(net299));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y0_300 (.LO(net300));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y0_301 (.LO(net301));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y15_302 (.LO(net302));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y15_303 (.LO(net303));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y15_304 (.LO(net304));
 sky130_fd_sc_hd__conb_1 arr_cell_x6_y15_305 (.LO(net305));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y0_306 (.LO(net306));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y0_307 (.LO(net307));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y0_308 (.LO(net308));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y15_309 (.LO(net309));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y15_310 (.LO(net310));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y15_311 (.LO(net311));
 sky130_fd_sc_hd__conb_1 arr_cell_x7_y15_312 (.LO(net312));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y0_313 (.LO(net313));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y0_314 (.LO(net314));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y0_315 (.LO(net315));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y15_316 (.LO(net316));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y15_317 (.LO(net317));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y15_318 (.LO(net318));
 sky130_fd_sc_hd__conb_1 arr_cell_x8_y15_319 (.LO(net319));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y0_320 (.LO(net320));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y0_321 (.LO(net321));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y0_322 (.LO(net322));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y15_323 (.LO(net323));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y15_324 (.LO(net324));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y15_325 (.LO(net325));
 sky130_fd_sc_hd__conb_1 arr_cell_x9_y15_326 (.LO(net326));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(reset),
    .X(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_08_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_13_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_13_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\cell_outs[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net56));
 sky130_ef_sc_hd__decap_12 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2472 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1913 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1916 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1928 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1940 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1561 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1817 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1830 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1861 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1872 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1901 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1905 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1914 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1918 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2169 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2173 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2219 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2231 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2257 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2517 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2537 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2601 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2685 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2699 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2711 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2729 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2737 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2993 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1264 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1432 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1612 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2134 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2300 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2129 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2297 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2305 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2489 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2509 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1959 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1981 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2005 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1761 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_2656 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_2834 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2984 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_2996 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2881 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_2885 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2891 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2896 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_2908 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1543 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1547 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_2421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_2431 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2447 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1517 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1521 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1535 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1545 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1683 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1713 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1717 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1721 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1725 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1729 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1755 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1785 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1809 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2349 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_2361 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2366 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2370 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2374 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2401 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2413 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2417 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2425 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_2429 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2431 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2443 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_2455 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_2656 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_2834 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1960 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_2133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1721 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1733 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1739 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1760 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2393 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_2405 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_2413 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2838 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2850 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_2862 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2996 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_2834 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_2838 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2842 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2848 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2860 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2884 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1761 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2433 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2437 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2996 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_2834 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_2838 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1960 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_2133 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1761 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1933 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1941 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_2101 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_2313 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_2483 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_2633 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2846 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2858 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1761 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2377 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_2381 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_2387 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_2391 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_2399 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_2403 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_2409 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2413 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_2781 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2981 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2993 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2999 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2846 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2858 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1397 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_2834 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_2838 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2996 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1761 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_2656 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_2834 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_290_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_292_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_292_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_297_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_299_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_299_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_300_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_302_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_304_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_306_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_306_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_306_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2838 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2850 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_2862 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_308_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2984 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_2996 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_310_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_314_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_318_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_320_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_320_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_320_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_1960 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_2133 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_320_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_322_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_324_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_324_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_326_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1721 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1733 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1739 ();
 sky130_fd_sc_hd__decap_4 FILLER_326_1760 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_2437 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_2445 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_330_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_333_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_333_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_334_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_2656 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_2834 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_340_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_340_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_346_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_349_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_350_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_352_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_355_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_357_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_357_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_359_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_360_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_2980 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_2992 ();
 sky130_fd_sc_hd__decap_4 FILLER_360_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_361_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_362_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_363_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_364_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_364_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_2656 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_2834 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_366_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_367_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_369_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_370_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_372_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_372_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_373_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_373_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_376_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_379_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_380_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_381_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_382_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_382_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_385_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_385_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_385_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_387_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_387_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_388_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1761 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_388_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_388_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_390_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_391_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_392_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_392_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2846 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2858 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_396_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_396_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_396_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_398_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_398_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_399_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_399_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_400_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_400_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_400_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_400_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_400_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_400_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_401_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_402_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_402_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_403_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_403_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_403_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_404_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_404_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_405_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_1960 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_2133 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_405_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_406_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_406_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_406_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_406_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_406_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_406_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_407_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_408_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_408_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_408_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_408_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_408_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_408_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_409_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_409_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_409_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_409_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_2968 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_2980 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_2988 ();
 sky130_fd_sc_hd__decap_4 FILLER_410_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_411_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_411_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_411_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_412_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_412_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_412_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_412_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_412_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_413_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_413_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_415_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_415_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_415_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_417_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_417_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_417_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_417_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_418_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_418_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_418_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_419_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_419_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_419_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_420_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_420_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_420_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_420_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_420_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_420_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_421_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_421_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_422_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_422_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_422_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_422_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_422_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_422_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_423_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_423_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_423_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_423_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_423_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_424_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_425_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_425_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_425_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_425_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_425_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2846 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2858 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_425_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_426_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_426_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_426_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_426_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_426_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_427_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_427_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_428_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_428_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_428_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_428_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_428_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_428_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_429_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_429_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_429_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_430_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_430_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_430_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_430_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_430_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_430_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_431_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_431_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_431_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_432_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_432_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_432_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_432_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2821 ();
 sky130_fd_sc_hd__decap_8 FILLER_432_2833 ();
 sky130_fd_sc_hd__fill_2 FILLER_432_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_432_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_433_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_433_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_433_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_434_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_434_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_434_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_434_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_434_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_435_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_435_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_435_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_435_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_435_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_435_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_435_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_436_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_436_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_437_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_437_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_437_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_437_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_437_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_438_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_438_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_439_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_439_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_439_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_440_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_440_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_440_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_440_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_440_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_440_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_441_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_441_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_441_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1761 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_1961 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2405 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_443_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_443_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_445_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_445_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_447_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_447_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_447_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_447_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_448_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_448_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_448_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_448_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_448_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_448_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_449_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_449_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_450_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_450_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_451_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_451_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_451_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_451_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_451_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_451_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_451_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_452_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_452_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_452_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_452_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_452_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_452_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_453_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_454_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_454_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_454_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_454_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_454_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_454_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_455_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_455_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_455_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_455_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_455_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_456_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_456_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_456_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_456_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_456_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_456_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_456_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_457_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_458_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_458_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_458_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_458_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_458_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_458_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_459_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_460_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_3010 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2821 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2833 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2845 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_462_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_462_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_462_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_462_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_462_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_463_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_463_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_463_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_463_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_463_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_463_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_463_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_464_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_464_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_464_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_464_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_464_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_464_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_465_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_465_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_465_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_465_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_465_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_465_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_465_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_466_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_466_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_467_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_467_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_467_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_468_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_468_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_468_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_468_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_468_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_468_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_469_2866 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_2870 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2872 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2884 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_2920 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_2926 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2928 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2940 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2952 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2964 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_2976 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_2982 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_2996 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_470_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_470_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_470_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_470_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_1600 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2122 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2296 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_470_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_2842 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2856 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2868 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_2892 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_2898 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2900 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2912 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2936 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_2948 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_2954 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2956 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2968 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2980 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_2992 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_3004 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_3010 ();
 sky130_fd_sc_hd__decap_4 FILLER_470_3012 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1536 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1545 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1557 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_1706 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1752 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1817 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1830 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1861 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_1872 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_1889 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1901 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1914 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_1926 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_1933 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1941 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2048 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2060 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2169 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2173 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2219 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_2231 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2253 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2257 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2313 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2414 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_2426 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2483 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2517 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2537 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2549 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2567 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2588 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2600 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2633 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2685 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2699 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2711 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2729 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2737 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2745 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_2757 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_2762 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_2770 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2101 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2135 ();
 sky130_fd_sc_hd__decap_8 FILLER_472_2147 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_473_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_473_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_473_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_475_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_475_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_475_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_477_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_477_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_477_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_478_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_478_1607 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_478_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_479_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_479_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_479_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_481_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_481_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_481_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_482_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_483_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_483_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_483_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_485_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_485_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_487_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_487_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_487_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_489_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_491_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_491_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_491_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_493_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_493_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_495_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_495_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_497_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_497_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_497_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_499_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_499_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_499_3013 ();
 sky130_fd_sc_hd__decap_8 FILLER_500_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_501_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_501_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_501_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_503_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_503_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_504_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_504_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_504_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2211 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_2221 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_3009 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_3015 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1331 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_2157 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2165 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2170 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2174 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2178 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2191 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2195 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2199 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2203 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2207 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2217 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2221 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2225 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_2229 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2741 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_2763 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_2997 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_3005 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_3008 ();
endmodule
