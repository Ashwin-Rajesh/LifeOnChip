VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO life_cell
  CLASS BLOCK ;
  FOREIGN life_cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 35.970 116.000 36.250 120.000 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END d
  PIN dl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END dl
  PIN dr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END dr
  PIN in_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END in_data
  PIN l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END l
  PIN load_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END load_in
  PIN load_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END load_out
  PIN out_data
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END out_data
  PIN prev_out_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 116.000 84.090 120.000 ;
    END
  END prev_out_data
  PIN r
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 58.520 120.000 59.120 ;
    END
  END r
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 104.760 120.000 105.360 ;
    END
  END reset
  PIN run
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 12.280 120.000 12.880 ;
    END
  END run
  PIN shift
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 35.400 120.000 36.000 ;
    END
  END shift
  PIN state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 81.640 120.000 82.240 ;
    END
  END state
  PIN u
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 116.000 60.170 120.000 ;
    END
  END u
  PIN ul
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.050 116.000 12.330 120.000 ;
    END
  END ul
  PIN ur
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.730 116.000 108.010 120.000 ;
    END
  END ur
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 4.670 10.640 114.080 109.040 ;
      LAYER met2 ;
        RECT 4.690 115.720 11.770 116.690 ;
        RECT 12.610 115.720 35.690 116.690 ;
        RECT 36.530 115.720 59.610 116.690 ;
        RECT 60.450 115.720 83.530 116.690 ;
        RECT 84.370 115.720 107.450 116.690 ;
        RECT 108.290 115.720 112.610 116.690 ;
        RECT 4.690 4.280 112.610 115.720 ;
        RECT 4.690 4.000 11.770 4.280 ;
        RECT 12.610 4.000 35.690 4.280 ;
        RECT 36.530 4.000 59.610 4.280 ;
        RECT 60.450 4.000 83.530 4.280 ;
        RECT 84.370 4.000 107.450 4.280 ;
        RECT 108.290 4.000 112.610 4.280 ;
      LAYER met3 ;
        RECT 4.000 105.760 116.000 108.965 ;
        RECT 4.400 104.360 115.600 105.760 ;
        RECT 4.000 82.640 116.000 104.360 ;
        RECT 4.400 81.240 115.600 82.640 ;
        RECT 4.000 59.520 116.000 81.240 ;
        RECT 4.400 58.120 115.600 59.520 ;
        RECT 4.000 36.400 116.000 58.120 ;
        RECT 4.400 35.000 115.600 36.400 ;
        RECT 4.000 13.280 116.000 35.000 ;
        RECT 4.400 11.880 115.600 13.280 ;
        RECT 4.000 10.715 116.000 11.880 ;
  END
END life_cell
END LIBRARY

