VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO life_cell
  CLASS BLOCK ;
  FOREIGN life_cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 40.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 27.220 10.640 28.820 27.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.720 10.640 16.320 27.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.720 10.640 41.320 27.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 15.270 36.000 15.550 40.000 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END d
  PIN dl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END dl
  PIN dr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END dr
  PIN in_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END in_data
  PIN l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END l
  PIN load_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END load_in
  PIN load_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END load_out
  PIN out_data
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END out_data
  PIN prev_out_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 34.590 36.000 34.870 40.000 ;
    END
  END prev_out_data
  PIN r
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 24.520 50.000 25.120 ;
    END
  END r
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 34.040 50.000 34.640 ;
    END
  END reset
  PIN run
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 5.480 50.000 6.080 ;
    END
  END run
  PIN shift
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 15.000 50.000 15.600 ;
    END
  END shift
  PIN state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END state
  PIN u
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 36.000 25.210 40.000 ;
    END
  END u
  PIN ul
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 5.610 36.000 5.890 40.000 ;
    END
  END ul
  PIN ur
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 36.000 44.530 40.000 ;
    END
  END ur
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 44.160 27.285 ;
      LAYER met1 ;
        RECT 4.670 10.640 44.550 27.440 ;
      LAYER met2 ;
        RECT 4.690 35.720 5.330 36.450 ;
        RECT 6.170 35.720 14.990 36.450 ;
        RECT 15.830 35.720 24.650 36.450 ;
        RECT 25.490 35.720 34.310 36.450 ;
        RECT 35.150 35.720 43.970 36.450 ;
        RECT 4.690 4.280 44.520 35.720 ;
        RECT 4.690 4.000 5.330 4.280 ;
        RECT 6.170 4.000 14.990 4.280 ;
        RECT 15.830 4.000 24.650 4.280 ;
        RECT 25.490 4.000 34.310 4.280 ;
        RECT 35.150 4.000 43.970 4.280 ;
      LAYER met3 ;
        RECT 4.400 33.640 45.600 34.505 ;
        RECT 4.000 25.520 46.000 33.640 ;
        RECT 4.400 24.120 45.600 25.520 ;
        RECT 4.000 16.000 46.000 24.120 ;
        RECT 4.400 14.600 45.600 16.000 ;
        RECT 4.000 6.480 46.000 14.600 ;
        RECT 4.400 5.615 45.600 6.480 ;
  END
END life_cell
END LIBRARY

